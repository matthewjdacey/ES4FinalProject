library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity jumbo is
        port (
                x : in unsigned(6 downto 0); -- 5bit for 32 pixel bird
                y : in unsigned(6 downto 0);
                rgb : out std_logic_vector(5 downto 0);
				clk : in std_logic
        );
end jumbo;

architecture synth of jumbo is
        signal smallx : unsigned(4 downto 0);
        signal smally : unsigned(4 downto 0);
begin
        smallx <= x(5 downto 1); -- divide to get image size (16x16)
        smally <= y(5 downto 1);

process(clk) begin
if rising_edge(clk) then
        rgb <=
			"000000" when smallx = "00000" and smally = "00000" else
			"000000" when smallx = "00001" and smally = "00000" else
			"000000" when smallx = "00010" and smally = "00000" else
			"000000" when smallx = "00011" and smally = "00000" else
			"000000" when smallx = "00100" and smally = "00000" else
			"000000" when smallx = "00101" and smally = "00000" else
			"000000" when smallx = "00110" and smally = "00000" else
			"000000" when smallx = "00111" and smally = "00000" else
			"000000" when smallx = "01000" and smally = "00000" else
			"000000" when smallx = "01001" and smally = "00000" else
			"000000" when smallx = "01010" and smally = "00000" else
			"000000" when smallx = "01011" and smally = "00000" else
			"000000" when smallx = "01100" and smally = "00000" else
			"000000" when smallx = "01101" and smally = "00000" else
			"000000" when smallx = "01110" and smally = "00000" else
			"000000" when smallx = "01111" and smally = "00000" else
			"000000" when smallx = "10000" and smally = "00000" else
			"000000" when smallx = "10001" and smally = "00000" else
			"000000" when smallx = "10010" and smally = "00000" else
			"000000" when smallx = "10011" and smally = "00000" else
			"000000" when smallx = "10100" and smally = "00000" else
			"000000" when smallx = "10101" and smally = "00000" else
			"000000" when smallx = "10110" and smally = "00000" else
			"000000" when smallx = "10111" and smally = "00000" else
			"000000" when smallx = "11000" and smally = "00000" else
			"000000" when smallx = "00000" and smally = "00001" else
			"000000" when smallx = "00001" and smally = "00001" else
			"000000" when smallx = "00010" and smally = "00001" else
			"000000" when smallx = "00011" and smally = "00001" else
			"000000" when smallx = "00100" and smally = "00001" else
			"000000" when smallx = "00101" and smally = "00001" else
			"000000" when smallx = "00110" and smally = "00001" else
			"000000" when smallx = "00111" and smally = "00001" else
			"000000" when smallx = "01000" and smally = "00001" else
			"000000" when smallx = "01001" and smally = "00001" else
			"000000" when smallx = "01010" and smally = "00001" else
			"000000" when smallx = "01011" and smally = "00001" else
			"000000" when smallx = "01100" and smally = "00001" else
			"000000" when smallx = "01101" and smally = "00001" else
			"000000" when smallx = "01110" and smally = "00001" else
			"000000" when smallx = "01111" and smally = "00001" else
			"000000" when smallx = "10000" and smally = "00001" else
			"000000" when smallx = "10001" and smally = "00001" else
			"000000" when smallx = "10010" and smally = "00001" else
			"000000" when smallx = "10011" and smally = "00001" else
			"000000" when smallx = "10100" and smally = "00001" else
			"000000" when smallx = "10101" and smally = "00001" else
			"000000" when smallx = "10110" and smally = "00001" else
			"000000" when smallx = "10111" and smally = "00001" else
			"000000" when smallx = "11000" and smally = "00001" else
			"000000" when smallx = "00000" and smally = "00010" else
			"000000" when smallx = "00001" and smally = "00010" else
			"000000" when smallx = "00010" and smally = "00010" else
			"000000" when smallx = "00011" and smally = "00010" else
			"000000" when smallx = "00100" and smally = "00010" else
			"000000" when smallx = "00101" and smally = "00010" else
			"000000" when smallx = "00110" and smally = "00010" else
			"000000" when smallx = "00111" and smally = "00010" else
			"000000" when smallx = "01000" and smally = "00010" else
			"000000" when smallx = "01001" and smally = "00010" else
			"000000" when smallx = "01010" and smally = "00010" else
			"000000" when smallx = "01011" and smally = "00010" else
			"000000" when smallx = "01100" and smally = "00010" else
			"000000" when smallx = "01101" and smally = "00010" else
			"000000" when smallx = "01110" and smally = "00010" else
			"000000" when smallx = "01111" and smally = "00010" else
			"000000" when smallx = "10000" and smally = "00010" else
			"000000" when smallx = "10001" and smally = "00010" else
			"000000" when smallx = "10010" and smally = "00010" else
			"000000" when smallx = "10011" and smally = "00010" else
			"000000" when smallx = "10100" and smally = "00010" else
			"000000" when smallx = "10101" and smally = "00010" else
			"000000" when smallx = "10110" and smally = "00010" else
			"000000" when smallx = "10111" and smally = "00010" else
			"000000" when smallx = "11000" and smally = "00010" else
			"000000" when smallx = "00000" and smally = "00011" else
			"000000" when smallx = "00001" and smally = "00011" else
			"000000" when smallx = "00010" and smally = "00011" else
			"000000" when smallx = "00011" and smally = "00011" else
			"000000" when smallx = "00100" and smally = "00011" else
			"000000" when smallx = "00101" and smally = "00011" else
			"000000" when smallx = "00110" and smally = "00011" else
			"000000" when smallx = "00111" and smally = "00011" else
			"000000" when smallx = "01000" and smally = "00011" else
			"000000" when smallx = "01001" and smally = "00011" else
			"000000" when smallx = "01010" and smally = "00011" else
			"000000" when smallx = "01011" and smally = "00011" else
			"000000" when smallx = "01100" and smally = "00011" else
			"000000" when smallx = "01101" and smally = "00011" else
			"000000" when smallx = "01110" and smally = "00011" else
			"000000" when smallx = "01111" and smally = "00011" else
			"000000" when smallx = "10000" and smally = "00011" else
			"000000" when smallx = "10001" and smally = "00011" else
			"000000" when smallx = "10010" and smally = "00011" else
			"000000" when smallx = "10011" and smally = "00011" else
			"000000" when smallx = "10100" and smally = "00011" else
			"000000" when smallx = "10101" and smally = "00011" else
			"000000" when smallx = "10110" and smally = "00011" else
			"000000" when smallx = "10111" and smally = "00011" else
			"000000" when smallx = "11000" and smally = "00011" else
			"000000" when smallx = "00000" and smally = "00100" else
			"000000" when smallx = "00001" and smally = "00100" else
			"000000" when smallx = "00010" and smally = "00100" else
			"000000" when smallx = "00011" and smally = "00100" else
			"000000" when smallx = "00100" and smally = "00100" else
			"000000" when smallx = "00101" and smally = "00100" else
			"000000" when smallx = "00110" and smally = "00100" else
			"000000" when smallx = "00111" and smally = "00100" else
			"000000" when smallx = "01000" and smally = "00100" else
			"000000" when smallx = "01001" and smally = "00100" else
			"000000" when smallx = "01010" and smally = "00100" else
			"000000" when smallx = "01011" and smally = "00100" else
			"000000" when smallx = "01100" and smally = "00100" else
			"000000" when smallx = "01101" and smally = "00100" else
			"000000" when smallx = "01110" and smally = "00100" else
			"000000" when smallx = "01111" and smally = "00100" else
			"000000" when smallx = "10000" and smally = "00100" else
			"000000" when smallx = "10001" and smally = "00100" else
			"000000" when smallx = "10010" and smally = "00100" else
			"000000" when smallx = "10011" and smally = "00100" else
			"000000" when smallx = "10100" and smally = "00100" else
			"000000" when smallx = "10101" and smally = "00100" else
			"000000" when smallx = "10110" and smally = "00100" else
			"000000" when smallx = "10111" and smally = "00100" else
			"000000" when smallx = "11000" and smally = "00100" else
			"000000" when smallx = "00000" and smally = "00101" else
			"000000" when smallx = "00001" and smally = "00101" else
			"000000" when smallx = "00010" and smally = "00101" else
			"000000" when smallx = "00011" and smally = "00101" else
			"000000" when smallx = "00100" and smally = "00101" else
			"000000" when smallx = "00101" and smally = "00101" else
			"000000" when smallx = "00110" and smally = "00101" else
			"000000" when smallx = "00111" and smally = "00101" else
			"000000" when smallx = "01000" and smally = "00101" else
			"101010" when smallx = "01001" and smally = "00101" else
			"101010" when smallx = "01010" and smally = "00101" else
			"101010" when smallx = "01011" and smally = "00101" else
			"101010" when smallx = "01100" and smally = "00101" else
			"101010" when smallx = "01101" and smally = "00101" else
			"101010" when smallx = "01110" and smally = "00101" else
			"101010" when smallx = "01111" and smally = "00101" else
			"101010" when smallx = "10000" and smally = "00101" else
			"101010" when smallx = "10001" and smally = "00101" else
			"101010" when smallx = "10010" and smally = "00101" else
			"000000" when smallx = "10011" and smally = "00101" else
			"000000" when smallx = "10100" and smally = "00101" else
			"000000" when smallx = "10101" and smally = "00101" else
			"000000" when smallx = "10110" and smally = "00101" else
			"000000" when smallx = "10111" and smally = "00101" else
			"000000" when smallx = "11000" and smally = "00101" else
			"000000" when smallx = "00000" and smally = "00110" else
			"000000" when smallx = "00001" and smally = "00110" else
			"000000" when smallx = "00010" and smally = "00110" else
			"000000" when smallx = "00011" and smally = "00110" else
			"000000" when smallx = "00100" and smally = "00110" else
			"000000" when smallx = "00101" and smally = "00110" else
			"101010" when smallx = "00110" and smally = "00110" else
			"101010" when smallx = "00111" and smally = "00110" else
			"101010" when smallx = "01000" and smally = "00110" else
			"010101" when smallx = "01001" and smally = "00110" else
			"010101" when smallx = "01010" and smally = "00110" else
			"010101" when smallx = "01011" and smally = "00110" else
			"010101" when smallx = "01100" and smally = "00110" else
			"010101" when smallx = "01101" and smally = "00110" else
			"010101" when smallx = "01110" and smally = "00110" else
			"010101" when smallx = "01111" and smally = "00110" else
			"101010" when smallx = "10000" and smally = "00110" else
			"101010" when smallx = "10001" and smally = "00110" else
			"101010" when smallx = "10010" and smally = "00110" else
			"101010" when smallx = "10011" and smally = "00110" else
			"000000" when smallx = "10100" and smally = "00110" else
			"000000" when smallx = "10101" and smally = "00110" else
			"000000" when smallx = "10110" and smally = "00110" else
			"000000" when smallx = "10111" and smally = "00110" else
			"000000" when smallx = "11000" and smally = "00110" else
			"000000" when smallx = "00000" and smally = "00111" else
			"000000" when smallx = "00001" and smally = "00111" else
			"000000" when smallx = "00010" and smally = "00111" else
			"000000" when smallx = "00011" and smally = "00111" else
			"000000" when smallx = "00100" and smally = "00111" else
			"000000" when smallx = "00101" and smally = "00111" else
			"101010" when smallx = "00110" and smally = "00111" else
			"101010" when smallx = "00111" and smally = "00111" else
			"010101" when smallx = "01000" and smally = "00111" else
			"010101" when smallx = "01001" and smally = "00111" else
			"010101" when smallx = "01010" and smally = "00111" else
			"010101" when smallx = "01011" and smally = "00111" else
			"010101" when smallx = "01100" and smally = "00111" else
			"010101" when smallx = "01101" and smally = "00111" else
			"010101" when smallx = "01110" and smally = "00111" else
			"010101" when smallx = "01111" and smally = "00111" else
			"101010" when smallx = "10000" and smally = "00111" else
			"101010" when smallx = "10001" and smally = "00111" else
			"101010" when smallx = "10010" and smally = "00111" else
			"101010" when smallx = "10011" and smally = "00111" else
			"000000" when smallx = "10100" and smally = "00111" else
			"000000" when smallx = "10101" and smally = "00111" else
			"000000" when smallx = "10110" and smally = "00111" else
			"000000" when smallx = "10111" and smally = "00111" else
			"000000" when smallx = "11000" and smally = "00111" else
			"000000" when smallx = "00000" and smally = "01000" else
			"000000" when smallx = "00001" and smally = "01000" else
			"000000" when smallx = "00010" and smally = "01000" else
			"101010" when smallx = "00011" and smally = "01000" else
			"101010" when smallx = "00100" and smally = "01000" else
			"101010" when smallx = "00101" and smally = "01000" else
			"101010" when smallx = "00110" and smally = "01000" else
			"101010" when smallx = "00111" and smally = "01000" else
			"010101" when smallx = "01000" and smally = "01000" else
			"010101" when smallx = "01001" and smally = "01000" else
			"010101" when smallx = "01010" and smally = "01000" else
			"010101" when smallx = "01011" and smally = "01000" else
			"010101" when smallx = "01100" and smally = "01000" else
			"010101" when smallx = "01101" and smally = "01000" else
			"101010" when smallx = "01110" and smally = "01000" else
			"101010" when smallx = "01111" and smally = "01000" else
			"101010" when smallx = "10000" and smally = "01000" else
			"101010" when smallx = "10001" and smally = "01000" else
			"101010" when smallx = "10010" and smally = "01000" else
			"101010" when smallx = "10011" and smally = "01000" else
			"000000" when smallx = "10100" and smally = "01000" else
			"000000" when smallx = "10101" and smally = "01000" else
			"000000" when smallx = "10110" and smally = "01000" else
			"000000" when smallx = "10111" and smally = "01000" else
			"000000" when smallx = "11000" and smally = "01000" else
			"000000" when smallx = "00000" and smally = "01001" else
			"000000" when smallx = "00001" and smally = "01001" else
			"000000" when smallx = "00010" and smally = "01001" else
			"101010" when smallx = "00011" and smally = "01001" else
			"101010" when smallx = "00100" and smally = "01001" else
			"101010" when smallx = "00101" and smally = "01001" else
			"101010" when smallx = "00110" and smally = "01001" else
			"101010" when smallx = "00111" and smally = "01001" else
			"010101" when smallx = "01000" and smally = "01001" else
			"010101" when smallx = "01001" and smally = "01001" else
			"010101" when smallx = "01010" and smally = "01001" else
			"010101" when smallx = "01011" and smally = "01001" else
			"010101" when smallx = "01100" and smally = "01001" else
			"010101" when smallx = "01101" and smally = "01001" else
			"101010" when smallx = "01110" and smally = "01001" else
			"101010" when smallx = "01111" and smally = "01001" else
			"101010" when smallx = "10000" and smally = "01001" else
			"101010" when smallx = "10001" and smally = "01001" else
			"101010" when smallx = "10010" and smally = "01001" else
			"101010" when smallx = "10011" and smally = "01001" else
			"000000" when smallx = "10100" and smally = "01001" else
			"000000" when smallx = "10101" and smally = "01001" else
			"000000" when smallx = "10110" and smally = "01001" else
			"000000" when smallx = "10111" and smally = "01001" else
			"000000" when smallx = "11000" and smally = "01001" else
			"000000" when smallx = "00000" and smally = "01010" else
			"000000" when smallx = "00001" and smally = "01010" else
			"000000" when smallx = "00010" and smally = "01010" else
			"101010" when smallx = "00011" and smally = "01010" else
			"101010" when smallx = "00100" and smally = "01010" else
			"101010" when smallx = "00101" and smally = "01010" else
			"101010" when smallx = "00110" and smally = "01010" else
			"101010" when smallx = "00111" and smally = "01010" else
			"010101" when smallx = "01000" and smally = "01010" else
			"010101" when smallx = "01001" and smally = "01010" else
			"010101" when smallx = "01010" and smally = "01010" else
			"010101" when smallx = "01011" and smally = "01010" else
			"010101" when smallx = "01100" and smally = "01010" else
			"010101" when smallx = "01101" and smally = "01010" else
			"101010" when smallx = "01110" and smally = "01010" else
			"101010" when smallx = "01111" and smally = "01010" else
			"101010" when smallx = "10000" and smally = "01010" else
			"101010" when smallx = "10001" and smally = "01010" else
			"101010" when smallx = "10010" and smally = "01010" else
			"101010" when smallx = "10011" and smally = "01010" else
			"000000" when smallx = "10100" and smally = "01010" else
			"000000" when smallx = "10101" and smally = "01010" else
			"000000" when smallx = "10110" and smally = "01010" else
			"000000" when smallx = "10111" and smally = "01010" else
			"000000" when smallx = "11000" and smally = "01010" else
			"000000" when smallx = "00000" and smally = "01011" else
			"000000" when smallx = "00001" and smally = "01011" else
			"101010" when smallx = "00010" and smally = "01011" else
			"101010" when smallx = "00011" and smally = "01011" else
			"101010" when smallx = "00100" and smally = "01011" else
			"101010" when smallx = "00101" and smally = "01011" else
			"101010" when smallx = "00110" and smally = "01011" else
			"101010" when smallx = "00111" and smally = "01011" else
			"101010" when smallx = "01000" and smally = "01011" else
			"101010" when smallx = "01001" and smally = "01011" else
			"101010" when smallx = "01010" and smally = "01011" else
			"101010" when smallx = "01011" and smally = "01011" else
			"101010" when smallx = "01100" and smally = "01011" else
			"101010" when smallx = "01101" and smally = "01011" else
			"101010" when smallx = "01110" and smally = "01011" else
			"101010" when smallx = "01111" and smally = "01011" else
			"010101" when smallx = "10000" and smally = "01011" else
			"101010" when smallx = "10001" and smally = "01011" else
			"101010" when smallx = "10010" and smally = "01011" else
			"101010" when smallx = "10011" and smally = "01011" else
			"000000" when smallx = "10100" and smally = "01011" else
			"000000" when smallx = "10101" and smally = "01011" else
			"000000" when smallx = "10110" and smally = "01011" else
			"000000" when smallx = "10111" and smally = "01011" else
			"000000" when smallx = "11000" and smally = "01011" else
			"101010" when smallx = "00000" and smally = "01100" else
			"101010" when smallx = "00001" and smally = "01100" else
			"101010" when smallx = "00010" and smally = "01100" else
			"101010" when smallx = "00011" and smally = "01100" else
			"101010" when smallx = "00100" and smally = "01100" else
			"101010" when smallx = "00101" and smally = "01100" else
			"101010" when smallx = "00110" and smally = "01100" else
			"101010" when smallx = "00111" and smally = "01100" else
			"101010" when smallx = "01000" and smally = "01100" else
			"101010" when smallx = "01001" and smally = "01100" else
			"101010" when smallx = "01010" and smally = "01100" else
			"101010" when smallx = "01011" and smally = "01100" else
			"101010" when smallx = "01100" and smally = "01100" else
			"101010" when smallx = "01101" and smally = "01100" else
			"101010" when smallx = "01110" and smally = "01100" else
			"101010" when smallx = "01111" and smally = "01100" else
			"101010" when smallx = "10000" and smally = "01100" else
			"101010" when smallx = "10001" and smally = "01100" else
			"101010" when smallx = "10010" and smally = "01100" else
			"101010" when smallx = "10011" and smally = "01100" else
			"000000" when smallx = "10100" and smally = "01100" else
			"000000" when smallx = "10101" and smally = "01100" else
			"000000" when smallx = "10110" and smally = "01100" else
			"000000" when smallx = "10111" and smally = "01100" else
			"000000" when smallx = "11000" and smally = "01100" else
			"101010" when smallx = "00000" and smally = "01101" else
			"101010" when smallx = "00001" and smally = "01101" else
			"101010" when smallx = "00010" and smally = "01101" else
			"101010" when smallx = "00011" and smally = "01101" else
			"101010" when smallx = "00100" and smally = "01101" else
			"101010" when smallx = "00101" and smally = "01101" else
			"101010" when smallx = "00110" and smally = "01101" else
			"101010" when smallx = "00111" and smally = "01101" else
			"101010" when smallx = "01000" and smally = "01101" else
			"101010" when smallx = "01001" and smally = "01101" else
			"101010" when smallx = "01010" and smally = "01101" else
			"101010" when smallx = "01011" and smally = "01101" else
			"101010" when smallx = "01100" and smally = "01101" else
			"101010" when smallx = "01101" and smally = "01101" else
			"101010" when smallx = "01110" and smally = "01101" else
			"101010" when smallx = "01111" and smally = "01101" else
			"101010" when smallx = "10000" and smally = "01101" else
			"101010" when smallx = "10001" and smally = "01101" else
			"101010" when smallx = "10010" and smally = "01101" else
			"101010" when smallx = "10011" and smally = "01101" else
			"000000" when smallx = "10100" and smally = "01101" else
			"000000" when smallx = "10101" and smally = "01101" else
			"101010" when smallx = "10110" and smally = "01101" else
			"000000" when smallx = "10111" and smally = "01101" else
			"000000" when smallx = "11000" and smally = "01101" else
			"000000" when smallx = "00000" and smally = "01110" else
			"000000" when smallx = "00001" and smally = "01110" else
			"101010" when smallx = "00010" and smally = "01110" else
			"101010" when smallx = "00011" and smally = "01110" else
			"101010" when smallx = "00100" and smally = "01110" else
			"101010" when smallx = "00101" and smally = "01110" else
			"101010" when smallx = "00110" and smally = "01110" else
			"101010" when smallx = "00111" and smally = "01110" else
			"101010" when smallx = "01000" and smally = "01110" else
			"101010" when smallx = "01001" and smally = "01110" else
			"101010" when smallx = "01010" and smally = "01110" else
			"101010" when smallx = "01011" and smally = "01110" else
			"101010" when smallx = "01100" and smally = "01110" else
			"101010" when smallx = "01101" and smally = "01110" else
			"101010" when smallx = "01110" and smally = "01110" else
			"101010" when smallx = "01111" and smally = "01110" else
			"101010" when smallx = "10000" and smally = "01110" else
			"101010" when smallx = "10001" and smally = "01110" else
			"101010" when smallx = "10010" and smally = "01110" else
			"101010" when smallx = "10011" and smally = "01110" else
			"000000" when smallx = "10100" and smally = "01110" else
			"101010" when smallx = "10101" and smally = "01110" else
			"101010" when smallx = "10110" and smally = "01110" else
			"101010" when smallx = "10111" and smally = "01110" else
			"000000" when smallx = "11000" and smally = "01110" else
			"000000" when smallx = "00000" and smally = "01111" else
			"000000" when smallx = "00001" and smally = "01111" else
			"101010" when smallx = "00010" and smally = "01111" else
			"101010" when smallx = "00011" and smally = "01111" else
			"101010" when smallx = "00100" and smally = "01111" else
			"101010" when smallx = "00101" and smally = "01111" else
			"101010" when smallx = "00110" and smally = "01111" else
			"101010" when smallx = "00111" and smally = "01111" else
			"101010" when smallx = "01000" and smally = "01111" else
			"101010" when smallx = "01001" and smally = "01111" else
			"101010" when smallx = "01010" and smally = "01111" else
			"101010" when smallx = "01011" and smally = "01111" else
			"101010" when smallx = "01100" and smally = "01111" else
			"101010" when smallx = "01101" and smally = "01111" else
			"101010" when smallx = "01110" and smally = "01111" else
			"101010" when smallx = "01111" and smally = "01111" else
			"101010" when smallx = "10000" and smally = "01111" else
			"101010" when smallx = "10001" and smally = "01111" else
			"101010" when smallx = "10010" and smally = "01111" else
			"101010" when smallx = "10011" and smally = "01111" else
			"101010" when smallx = "10100" and smally = "01111" else
			"101010" when smallx = "10101" and smally = "01111" else
			"101010" when smallx = "10110" and smally = "01111" else
			"000000" when smallx = "10111" and smally = "01111" else
			"000000" when smallx = "11000" and smally = "01111" else
			"000000" when smallx = "00000" and smally = "10000" else
			"000000" when smallx = "00001" and smally = "10000" else
			"101010" when smallx = "00010" and smally = "10000" else
			"101010" when smallx = "00011" and smally = "10000" else
			"101010" when smallx = "00100" and smally = "10000" else
			"101010" when smallx = "00101" and smally = "10000" else
			"101010" when smallx = "00110" and smally = "10000" else
			"101010" when smallx = "00111" and smally = "10000" else
			"101010" when smallx = "01000" and smally = "10000" else
			"101010" when smallx = "01001" and smally = "10000" else
			"101010" when smallx = "01010" and smally = "10000" else
			"101010" when smallx = "01011" and smally = "10000" else
			"101010" when smallx = "01100" and smally = "10000" else
			"101010" when smallx = "01101" and smally = "10000" else
			"101010" when smallx = "01110" and smally = "10000" else
			"101010" when smallx = "01111" and smally = "10000" else
			"101010" when smallx = "10000" and smally = "10000" else
			"101010" when smallx = "10001" and smally = "10000" else
			"101010" when smallx = "10010" and smally = "10000" else
			"101010" when smallx = "10011" and smally = "10000" else
			"101010" when smallx = "10100" and smally = "10000" else
			"101010" when smallx = "10101" and smally = "10000" else
			"000000" when smallx = "10110" and smally = "10000" else
			"000000" when smallx = "10111" and smally = "10000" else
			"000000" when smallx = "11000" and smally = "10000" else
			"000000" when smallx = "00000" and smally = "10001" else
			"000000" when smallx = "00001" and smally = "10001" else
			"101010" when smallx = "00010" and smally = "10001" else
			"101010" when smallx = "00011" and smally = "10001" else
			"101010" when smallx = "00100" and smally = "10001" else
			"101010" when smallx = "00101" and smally = "10001" else
			"101010" when smallx = "00110" and smally = "10001" else
			"101010" when smallx = "00111" and smally = "10001" else
			"000000" when smallx = "01000" and smally = "10001" else
			"000000" when smallx = "01001" and smally = "10001" else
			"000000" when smallx = "01010" and smally = "10001" else
			"101010" when smallx = "01011" and smally = "10001" else
			"101010" when smallx = "01100" and smally = "10001" else
			"101010" when smallx = "01101" and smally = "10001" else
			"101010" when smallx = "01110" and smally = "10001" else
			"101010" when smallx = "01111" and smally = "10001" else
			"101010" when smallx = "10000" and smally = "10001" else
			"000000" when smallx = "10001" and smally = "10001" else
			"000000" when smallx = "10010" and smally = "10001" else
			"000000" when smallx = "10011" and smally = "10001" else
			"000000" when smallx = "10100" and smally = "10001" else
			"000000" when smallx = "10101" and smally = "10001" else
			"000000" when smallx = "10110" and smally = "10001" else
			"000000" when smallx = "10111" and smally = "10001" else
			"000000" when smallx = "11000" and smally = "10001" else
			"000000" when smallx = "00000" and smally = "10010" else
			"000000" when smallx = "00001" and smally = "10010" else
			"101010" when smallx = "00010" and smally = "10010" else
			"101010" when smallx = "00011" and smally = "10010" else
			"101010" when smallx = "00100" and smally = "10010" else
			"101010" when smallx = "00101" and smally = "10010" else
			"101010" when smallx = "00110" and smally = "10010" else
			"101010" when smallx = "00111" and smally = "10010" else
			"000000" when smallx = "01000" and smally = "10010" else
			"000000" when smallx = "01001" and smally = "10010" else
			"000000" when smallx = "01010" and smally = "10010" else
			"101010" when smallx = "01011" and smally = "10010" else
			"101010" when smallx = "01100" and smally = "10010" else
			"101010" when smallx = "01101" and smally = "10010" else
			"101010" when smallx = "01110" and smally = "10010" else
			"101010" when smallx = "01111" and smally = "10010" else
			"101010" when smallx = "10000" and smally = "10010" else
			"000000" when smallx = "10001" and smally = "10010" else
			"000000" when smallx = "10010" and smally = "10010" else
			"000000" when smallx = "10011" and smally = "10010" else
			"000000" when smallx = "10100" and smally = "10010" else
			"000000" when smallx = "10101" and smally = "10010" else
			"000000" when smallx = "10110" and smally = "10010" else
			"000000" when smallx = "10111" and smally = "10010" else
			"000000" when smallx = "11000" and smally = "10010" else
			"000000" when smallx = "00000" and smally = "10011" else
			"000000" when smallx = "00001" and smally = "10011" else
			"101010" when smallx = "00010" and smally = "10011" else
			"101010" when smallx = "00011" and smally = "10011" else
			"101010" when smallx = "00100" and smally = "10011" else
			"101010" when smallx = "00101" and smally = "10011" else
			"101010" when smallx = "00110" and smally = "10011" else
			"101010" when smallx = "00111" and smally = "10011" else
			"000000" when smallx = "01000" and smally = "10011" else
			"000000" when smallx = "01001" and smally = "10011" else
			"000000" when smallx = "01010" and smally = "10011" else
			"101010" when smallx = "01011" and smally = "10011" else
			"101010" when smallx = "01100" and smally = "10011" else
			"101010" when smallx = "01101" and smally = "10011" else
			"101010" when smallx = "01110" and smally = "10011" else
			"101010" when smallx = "01111" and smally = "10011" else
			"101010" when smallx = "10000" and smally = "10011" else
			"000000" when smallx = "10001" and smally = "10011" else
			"000000" when smallx = "10010" and smally = "10011" else
			"000000" when smallx = "10011" and smally = "10011" else
			"000000" when smallx = "10100" and smally = "10011" else
			"000000" when smallx = "10101" and smally = "10011" else
			"000000" when smallx = "10110" and smally = "10011" else
			"000000" when smallx = "10111" and smally = "10011" else
			"000000" when smallx = "11000" and smally = "10011" else
			"000000" when smallx = "00000" and smally = "10100" else
			"000000" when smallx = "00001" and smally = "10100" else
			"101010" when smallx = "00010" and smally = "10100" else
			"101010" when smallx = "00011" and smally = "10100" else
			"101010" when smallx = "00100" and smally = "10100" else
			"101010" when smallx = "00101" and smally = "10100" else
			"101010" when smallx = "00110" and smally = "10100" else
			"101010" when smallx = "00111" and smally = "10100" else
			"000000" when smallx = "01000" and smally = "10100" else
			"000000" when smallx = "01001" and smally = "10100" else
			"000000" when smallx = "01010" and smally = "10100" else
			"101010" when smallx = "01011" and smally = "10100" else
			"101010" when smallx = "01100" and smally = "10100" else
			"101010" when smallx = "01101" and smally = "10100" else
			"101010" when smallx = "01110" and smally = "10100" else
			"101010" when smallx = "01111" and smally = "10100" else
			"101010" when smallx = "10000" and smally = "10100" else
			"000000" when smallx = "10001" and smally = "10100" else
			"000000" when smallx = "10010" and smally = "10100" else
			"000000" when smallx = "10011" and smally = "10100" else
			"000000" when smallx = "10100" and smally = "10100" else
			"000000" when smallx = "10101" and smally = "10100" else
			"000000" when smallx = "10110" and smally = "10100" else
			"000000" when smallx = "10111" and smally = "10100" else
			"000000" when smallx = "11000" and smally = "10100" else
			"000000" when smallx = "00000" and smally = "10101" else
			"000000" when smallx = "00001" and smally = "10101" else
			"101010" when smallx = "00010" and smally = "10101" else
			"101010" when smallx = "00011" and smally = "10101" else
			"101010" when smallx = "00100" and smally = "10101" else
			"101010" when smallx = "00101" and smally = "10101" else
			"101010" when smallx = "00110" and smally = "10101" else
			"101010" when smallx = "00111" and smally = "10101" else
			"000000" when smallx = "01000" and smally = "10101" else
			"000000" when smallx = "01001" and smally = "10101" else
			"000000" when smallx = "01010" and smally = "10101" else
			"101010" when smallx = "01011" and smally = "10101" else
			"101010" when smallx = "01100" and smally = "10101" else
			"101010" when smallx = "01101" and smally = "10101" else
			"101010" when smallx = "01110" and smally = "10101" else
			"101010" when smallx = "01111" and smally = "10101" else
			"101010" when smallx = "10000" and smally = "10101" else
			"000000" when smallx = "10001" and smally = "10101" else
			"000000" when smallx = "10010" and smally = "10101" else
			"000000" when smallx = "10011" and smally = "10101" else
			"000000" when smallx = "10100" and smally = "10101" else
			"000000" when smallx = "10101" and smally = "10101" else
			"000000" when smallx = "10110" and smally = "10101" else
			"000000" when smallx = "10111" and smally = "10101" else
			"000000" when smallx = "11000" and smally = "10101" else
			"000000" when smallx = "00000" and smally = "10110" else
			"000000" when smallx = "00001" and smally = "10110" else
			"000000" when smallx = "00010" and smally = "10110" else
			"000000" when smallx = "00011" and smally = "10110" else
			"000000" when smallx = "00100" and smally = "10110" else
			"000000" when smallx = "00101" and smally = "10110" else
			"000000" when smallx = "00110" and smally = "10110" else
			"000000" when smallx = "00111" and smally = "10110" else
			"000000" when smallx = "01000" and smally = "10110" else
			"000000" when smallx = "01001" and smally = "10110" else
			"000000" when smallx = "01010" and smally = "10110" else
			"000000" when smallx = "01011" and smally = "10110" else
			"000000" when smallx = "01100" and smally = "10110" else
			"000000" when smallx = "01101" and smally = "10110" else
			"000000" when smallx = "01110" and smally = "10110" else
			"000000" when smallx = "01111" and smally = "10110" else
			"000000" when smallx = "10000" and smally = "10110" else
			"000000" when smallx = "10001" and smally = "10110" else
			"000000" when smallx = "10010" and smally = "10110" else
			"000000" when smallx = "10011" and smally = "10110" else
			"000000" when smallx = "10100" and smally = "10110" else
			"000000" when smallx = "10101" and smally = "10110" else
			"000000" when smallx = "10110" and smally = "10110" else
			"000000" when smallx = "10111" and smally = "10110" else
			"000000" when smallx = "11000" and smally = "10110" else
			"000000" when smallx = "00000" and smally = "10111" else
			"000000" when smallx = "00001" and smally = "10111" else
			"000000" when smallx = "00010" and smally = "10111" else
			"000000" when smallx = "00011" and smally = "10111" else
			"000000" when smallx = "00100" and smally = "10111" else
			"000000" when smallx = "00101" and smally = "10111" else
			"000000" when smallx = "00110" and smally = "10111" else
			"000000" when smallx = "00111" and smally = "10111" else
			"000000" when smallx = "01000" and smally = "10111" else
			"000000" when smallx = "01001" and smally = "10111" else
			"000000" when smallx = "01010" and smally = "10111" else
			"000000" when smallx = "01011" and smally = "10111" else
			"000000" when smallx = "01100" and smally = "10111" else
			"000000" when smallx = "01101" and smally = "10111" else
			"000000" when smallx = "01110" and smally = "10111" else
			"000000" when smallx = "01111" and smally = "10111" else
			"000000" when smallx = "10000" and smally = "10111" else
			"000000" when smallx = "10001" and smally = "10111" else
			"000000" when smallx = "10010" and smally = "10111" else
			"000000" when smallx = "10011" and smally = "10111" else
			"000000" when smallx = "10100" and smally = "10111" else
			"000000" when smallx = "10101" and smally = "10111" else
			"000000" when smallx = "10110" and smally = "10111" else
			"000000" when smallx = "10111" and smally = "10111" else
			"000000" when smallx = "11000" and smally = "10111" else
			"000000" when smallx = "00000" and smally = "11000" else
			"000000" when smallx = "00001" and smally = "11000" else
			"000000" when smallx = "00010" and smally = "11000" else
			"000000" when smallx = "00011" and smally = "11000" else
			"000000" when smallx = "00100" and smally = "11000" else
			"000000" when smallx = "00101" and smally = "11000" else
			"000000" when smallx = "00110" and smally = "11000" else
			"000000" when smallx = "00111" and smally = "11000" else
			"000000" when smallx = "01000" and smally = "11000" else
			"000000" when smallx = "01001" and smally = "11000" else
			"000000" when smallx = "01010" and smally = "11000" else
			"000000" when smallx = "01011" and smally = "11000" else
			"000000" when smallx = "01100" and smally = "11000" else
			"000000" when smallx = "01101" and smally = "11000" else
			"000000" when smallx = "01110" and smally = "11000" else
			"000000" when smallx = "01111" and smally = "11000" else
			"000000" when smallx = "10000" and smally = "11000" else
			"000000" when smallx = "10001" and smally = "11000" else
			"000000" when smallx = "10010" and smally = "11000" else
			"000000" when smallx = "10011" and smally = "11000" else
			"000000" when smallx = "10100" and smally = "11000" else
			"000000" when smallx = "10101" and smally = "11000" else
			"000000" when smallx = "10110" and smally = "11000" else
			"000000" when smallx = "10111" and smally = "11000" else
			"000000" when smallx = "11000" and smally = "11000" else
			"000011";
end if;
end process;
end;
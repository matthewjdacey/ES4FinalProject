library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity jumbo is
        port (
                x : in unsigned(9 downto 0); -- 5bit for 32 pixel bird
                y : in unsigned(9 downto 0);
                rgb : out std_logic_vector(5 downto 0);
				clk : in std_logic
        );
end jumbo;

architecture synth of jumbo is
        signal smallx : unsigned(7 downto 0);
        signal smally : unsigned(7 downto 0);
begin
        smallx <= x(8 downto 1); -- divide to get image size (16x16)
        smally <= y(8 downto 1);

process(clk) begin
if rising_edge(clk) then
        rgb <=
			"011011" when smallx = "0000000" and smally = "0000000" else
			"011011" when smallx = "0000001" and smally = "0000000" else
			"011011" when smallx = "0000010" and smally = "0000000" else
			"011011" when smallx = "0000011" and smally = "0000000" else
			"011011" when smallx = "0000100" and smally = "0000000" else
			"011011" when smallx = "0000101" and smally = "0000000" else
			"011011" when smallx = "0000110" and smally = "0000000" else
			"011011" when smallx = "0000111" and smally = "0000000" else
			"000000" when smallx = "0001000" and smally = "0000000" else
			"000000" when smallx = "0001001" and smally = "0000000" else
			"000000" when smallx = "0001010" and smally = "0000000" else
			"000000" when smallx = "0001011" and smally = "0000000" else
			"000000" when smallx = "0001100" and smally = "0000000" else
			"000000" when smallx = "0001101" and smally = "0000000" else
			"000000" when smallx = "0001110" and smally = "0000000" else
			"000000" when smallx = "0001111" and smally = "0000000" else
			"011011" when smallx = "0010000" and smally = "0000000" else
			"011011" when smallx = "0010001" and smally = "0000000" else
			"011011" when smallx = "0010010" and smally = "0000000" else
			"011011" when smallx = "0010011" and smally = "0000000" else
			"011011" when smallx = "0010100" and smally = "0000000" else
			"011011" when smallx = "0010101" and smally = "0000000" else
			"011011" when smallx = "0000000" and smally = "0000001" else
			"011011" when smallx = "0000001" and smally = "0000001" else
			"011011" when smallx = "0000010" and smally = "0000001" else
			"011011" when smallx = "0000011" and smally = "0000001" else
			"011011" when smallx = "0000100" and smally = "0000001" else
			"011011" when smallx = "0000101" and smally = "0000001" else
			"011011" when smallx = "0000110" and smally = "0000001" else
			"000000" when smallx = "0000111" and smally = "0000001" else
			"010101" when smallx = "0001000" and smally = "0000001" else
			"010101" when smallx = "0001001" and smally = "0000001" else
			"010101" when smallx = "0001010" and smally = "0000001" else
			"010101" when smallx = "0001011" and smally = "0000001" else
			"010101" when smallx = "0001100" and smally = "0000001" else
			"000000" when smallx = "0001101" and smally = "0000001" else
			"101010" when smallx = "0001110" and smally = "0000001" else
			"101010" when smallx = "0001111" and smally = "0000001" else
			"000000" when smallx = "0010000" and smally = "0000001" else
			"011011" when smallx = "0010001" and smally = "0000001" else
			"011011" when smallx = "0010010" and smally = "0000001" else
			"011011" when smallx = "0010011" and smally = "0000001" else
			"011011" when smallx = "0010100" and smally = "0000001" else
			"011011" when smallx = "0010101" and smally = "0000001" else
			"011011" when smallx = "0000000" and smally = "0000010" else
			"011011" when smallx = "0000001" and smally = "0000010" else
			"011011" when smallx = "0000010" and smally = "0000010" else
			"011011" when smallx = "0000011" and smally = "0000010" else
			"000000" when smallx = "0000100" and smally = "0000010" else
			"000000" when smallx = "0000101" and smally = "0000010" else
			"000000" when smallx = "0000110" and smally = "0000010" else
			"000000" when smallx = "0000111" and smally = "0000010" else
			"010101" when smallx = "0001000" and smally = "0000010" else
			"010101" when smallx = "0001001" and smally = "0000010" else
			"010101" when smallx = "0001010" and smally = "0000010" else
			"010101" when smallx = "0001011" and smally = "0000010" else
			"010101" when smallx = "0001100" and smally = "0000010" else
			"000000" when smallx = "0001101" and smally = "0000010" else
			"101010" when smallx = "0001110" and smally = "0000010" else
			"101010" when smallx = "0001111" and smally = "0000010" else
			"101010" when smallx = "0010000" and smally = "0000010" else
			"000000" when smallx = "0010001" and smally = "0000010" else
			"011011" when smallx = "0010010" and smally = "0000010" else
			"011011" when smallx = "0010011" and smally = "0000010" else
			"011011" when smallx = "0010100" and smally = "0000010" else
			"011011" when smallx = "0010101" and smally = "0000010" else
			"011011" when smallx = "0000000" and smally = "0000011" else
			"011011" when smallx = "0000001" and smally = "0000011" else
			"011011" when smallx = "0000010" and smally = "0000011" else
			"000000" when smallx = "0000011" and smally = "0000011" else
			"101010" when smallx = "0000100" and smally = "0000011" else
			"101010" when smallx = "0000101" and smally = "0000011" else
			"101010" when smallx = "0000110" and smally = "0000011" else
			"101010" when smallx = "0000111" and smally = "0000011" else
			"000000" when smallx = "0001000" and smally = "0000011" else
			"010101" when smallx = "0001001" and smally = "0000011" else
			"010101" when smallx = "0001010" and smally = "0000011" else
			"010101" when smallx = "0001011" and smally = "0000011" else
			"000000" when smallx = "0001100" and smally = "0000011" else
			"101010" when smallx = "0001101" and smally = "0000011" else
			"101010" when smallx = "0001110" and smally = "0000011" else
			"101010" when smallx = "0001111" and smally = "0000011" else
			"101010" when smallx = "0010000" and smally = "0000011" else
			"000000" when smallx = "0010001" and smally = "0000011" else
			"011011" when smallx = "0010010" and smally = "0000011" else
			"011011" when smallx = "0010011" and smally = "0000011" else
			"011011" when smallx = "0010100" and smally = "0000011" else
			"011011" when smallx = "0010101" and smally = "0000011" else
			"011011" when smallx = "0000000" and smally = "0000100" else
			"011011" when smallx = "0000001" and smally = "0000100" else
			"000000" when smallx = "0000010" and smally = "0000100" else
			"101010" when smallx = "0000011" and smally = "0000100" else
			"101010" when smallx = "0000100" and smally = "0000100" else
			"101010" when smallx = "0000101" and smally = "0000100" else
			"101010" when smallx = "0000110" and smally = "0000100" else
			"101010" when smallx = "0000111" and smally = "0000100" else
			"101010" when smallx = "0001000" and smally = "0000100" else
			"000000" when smallx = "0001001" and smally = "0000100" else
			"000000" when smallx = "0001010" and smally = "0000100" else
			"000000" when smallx = "0001011" and smally = "0000100" else
			"101010" when smallx = "0001100" and smally = "0000100" else
			"101010" when smallx = "0001101" and smally = "0000100" else
			"101010" when smallx = "0001110" and smally = "0000100" else
			"101010" when smallx = "0001111" and smally = "0000100" else
			"101010" when smallx = "0010000" and smally = "0000100" else
			"000000" when smallx = "0010001" and smally = "0000100" else
			"011011" when smallx = "0010010" and smally = "0000100" else
			"011011" when smallx = "0010011" and smally = "0000100" else
			"011011" when smallx = "0010100" and smally = "0000100" else
			"011011" when smallx = "0010101" and smally = "0000100" else
			"011011" when smallx = "0000000" and smally = "0000101" else
			"011011" when smallx = "0000001" and smally = "0000101" else
			"000000" when smallx = "0000010" and smally = "0000101" else
			"101010" when smallx = "0000011" and smally = "0000101" else
			"101010" when smallx = "0000100" and smally = "0000101" else
			"101010" when smallx = "0000101" and smally = "0000101" else
			"101010" when smallx = "0000110" and smally = "0000101" else
			"101010" when smallx = "0000111" and smally = "0000101" else
			"101010" when smallx = "0001000" and smally = "0000101" else
			"101010" when smallx = "0001001" and smally = "0000101" else
			"101010" when smallx = "0001010" and smally = "0000101" else
			"101010" when smallx = "0001011" and smally = "0000101" else
			"101010" when smallx = "0001100" and smally = "0000101" else
			"101010" when smallx = "0001101" and smally = "0000101" else
			"101010" when smallx = "0001110" and smally = "0000101" else
			"000000" when smallx = "0001111" and smally = "0000101" else
			"101010" when smallx = "0010000" and smally = "0000101" else
			"000000" when smallx = "0010001" and smally = "0000101" else
			"011011" when smallx = "0010010" and smally = "0000101" else
			"000000" when smallx = "0010011" and smally = "0000101" else
			"000000" when smallx = "0010100" and smally = "0000101" else
			"011011" when smallx = "0010101" and smally = "0000101" else
			"000000" when smallx = "0000000" and smally = "0000110" else
			"000000" when smallx = "0000001" and smally = "0000110" else
			"000000" when smallx = "0000010" and smally = "0000110" else
			"101010" when smallx = "0000011" and smally = "0000110" else
			"101010" when smallx = "0000100" and smally = "0000110" else
			"101010" when smallx = "0000101" and smally = "0000110" else
			"101010" when smallx = "0000110" and smally = "0000110" else
			"101010" when smallx = "0000111" and smally = "0000110" else
			"101010" when smallx = "0001000" and smally = "0000110" else
			"101010" when smallx = "0001001" and smally = "0000110" else
			"101010" when smallx = "0001010" and smally = "0000110" else
			"101010" when smallx = "0001011" and smally = "0000110" else
			"101010" when smallx = "0001100" and smally = "0000110" else
			"101010" when smallx = "0001101" and smally = "0000110" else
			"101010" when smallx = "0001110" and smally = "0000110" else
			"101010" when smallx = "0001111" and smally = "0000110" else
			"101010" when smallx = "0010000" and smally = "0000110" else
			"000000" when smallx = "0010001" and smally = "0000110" else
			"000000" when smallx = "0010010" and smally = "0000110" else
			"101010" when smallx = "0010011" and smally = "0000110" else
			"101010" when smallx = "0010100" and smally = "0000110" else
			"000000" when smallx = "0010101" and smally = "0000110" else
			"011011" when smallx = "0000000" and smally = "0000111" else
			"011011" when smallx = "0000001" and smally = "0000111" else
			"000000" when smallx = "0000010" and smally = "0000111" else
			"101010" when smallx = "0000011" and smally = "0000111" else
			"101010" when smallx = "0000100" and smally = "0000111" else
			"101010" when smallx = "0000101" and smally = "0000111" else
			"101010" when smallx = "0000110" and smally = "0000111" else
			"101010" when smallx = "0000111" and smally = "0000111" else
			"101010" when smallx = "0001000" and smally = "0000111" else
			"101010" when smallx = "0001001" and smally = "0000111" else
			"101010" when smallx = "0001010" and smally = "0000111" else
			"101010" when smallx = "0001011" and smally = "0000111" else
			"101010" when smallx = "0001100" and smally = "0000111" else
			"101010" when smallx = "0001101" and smally = "0000111" else
			"101010" when smallx = "0001110" and smally = "0000111" else
			"101010" when smallx = "0001111" and smally = "0000111" else
			"101010" when smallx = "0010000" and smally = "0000111" else
			"101010" when smallx = "0010001" and smally = "0000111" else
			"101010" when smallx = "0010010" and smally = "0000111" else
			"101010" when smallx = "0010011" and smally = "0000111" else
			"000000" when smallx = "0010100" and smally = "0000111" else
			"011011" when smallx = "0010101" and smally = "0000111" else
			"011011" when smallx = "0000000" and smally = "0001000" else
			"011011" when smallx = "0000001" and smally = "0001000" else
			"000000" when smallx = "0000010" and smally = "0001000" else
			"101010" when smallx = "0000011" and smally = "0001000" else
			"101010" when smallx = "0000100" and smally = "0001000" else
			"000000" when smallx = "0000101" and smally = "0001000" else
			"000000" when smallx = "0000110" and smally = "0001000" else
			"000000" when smallx = "0000111" and smally = "0001000" else
			"000000" when smallx = "0001000" and smally = "0001000" else
			"000000" when smallx = "0001001" and smally = "0001000" else
			"000000" when smallx = "0001010" and smally = "0001000" else
			"000000" when smallx = "0001011" and smally = "0001000" else
			"101010" when smallx = "0001100" and smally = "0001000" else
			"101010" when smallx = "0001101" and smally = "0001000" else
			"101010" when smallx = "0001110" and smally = "0001000" else
			"101010" when smallx = "0001111" and smally = "0001000" else
			"101010" when smallx = "0010000" and smally = "0001000" else
			"000000" when smallx = "0010001" and smally = "0001000" else
			"000000" when smallx = "0010010" and smally = "0001000" else
			"000000" when smallx = "0010011" and smally = "0001000" else
			"011011" when smallx = "0010100" and smally = "0001000" else
			"011011" when smallx = "0010101" and smally = "0001000" else
			"011011" when smallx = "0000000" and smally = "0001001" else
			"011011" when smallx = "0000001" and smally = "0001001" else
			"000000" when smallx = "0000010" and smally = "0001001" else
			"101010" when smallx = "0000011" and smally = "0001001" else
			"101010" when smallx = "0000100" and smally = "0001001" else
			"000000" when smallx = "0000101" and smally = "0001001" else
			"011011" when smallx = "0000110" and smally = "0001001" else
			"011011" when smallx = "0000111" and smally = "0001001" else
			"011011" when smallx = "0001000" and smally = "0001001" else
			"011011" when smallx = "0001001" and smally = "0001001" else
			"011011" when smallx = "0001010" and smally = "0001001" else
			"000000" when smallx = "0001011" and smally = "0001001" else
			"101010" when smallx = "0001100" and smally = "0001001" else
			"101010" when smallx = "0001101" and smally = "0001001" else
			"000000" when smallx = "0001110" and smally = "0001001" else
			"000000" when smallx = "0001111" and smally = "0001001" else
			"000000" when smallx = "0010000" and smally = "0001001" else
			"011011" when smallx = "0010001" and smally = "0001001" else
			"011011" when smallx = "0010010" and smally = "0001001" else
			"011011" when smallx = "0010011" and smally = "0001001" else
			"011011" when smallx = "0010100" and smally = "0001001" else
			"011011" when smallx = "0010101" and smally = "0001001" else
			"011011" when smallx = "0000000" and smally = "0001010" else
			"011011" when smallx = "0000001" and smally = "0001010" else
			"000000" when smallx = "0000010" and smally = "0001010" else
			"101010" when smallx = "0000011" and smally = "0001010" else
			"101010" when smallx = "0000100" and smally = "0001010" else
			"000000" when smallx = "0000101" and smally = "0001010" else
			"011011" when smallx = "0000110" and smally = "0001010" else
			"011011" when smallx = "0000111" and smally = "0001010" else
			"011011" when smallx = "0001000" and smally = "0001010" else
			"011011" when smallx = "0001001" and smally = "0001010" else
			"011011" when smallx = "0001010" and smally = "0001010" else
			"000000" when smallx = "0001011" and smally = "0001010" else
			"101010" when smallx = "0001100" and smally = "0001010" else
			"101010" when smallx = "0001101" and smally = "0001010" else
			"000000" when smallx = "0001110" and smally = "0001010" else
			"011011" when smallx = "0001111" and smally = "0001010" else
			"011011" when smallx = "0010000" and smally = "0001010" else
			"011011" when smallx = "0010001" and smally = "0001010" else
			"011011" when smallx = "0010010" and smally = "0001010" else
			"011011" when smallx = "0010011" and smally = "0001010" else
			"011011" when smallx = "0010100" and smally = "0001010" else
			"011011" when smallx = "0010101" and smally = "0001010" else
			"011011" when smallx = "0000000" and smally = "0001011" else
			"011011" when smallx = "0000001" and smally = "0001011" else
			"000000" when smallx = "0000010" and smally = "0001011" else
			"101010" when smallx = "0000011" and smally = "0001011" else
			"101010" when smallx = "0000100" and smally = "0001011" else
			"000000" when smallx = "0000101" and smally = "0001011" else
			"011011" when smallx = "0000110" and smally = "0001011" else
			"011011" when smallx = "0000111" and smally = "0001011" else
			"011011" when smallx = "0001000" and smally = "0001011" else
			"011011" when smallx = "0001001" and smally = "0001011" else
			"011011" when smallx = "0001010" and smally = "0001011" else
			"000000" when smallx = "0001011" and smally = "0001011" else
			"101010" when smallx = "0001100" and smally = "0001011" else
			"101010" when smallx = "0001101" and smally = "0001011" else
			"000000" when smallx = "0001110" and smally = "0001011" else
			"011011" when smallx = "0001111" and smally = "0001011" else
			"011011" when smallx = "0010000" and smally = "0001011" else
			"011011" when smallx = "0010001" and smally = "0001011" else
			"011011" when smallx = "0010010" and smally = "0001011" else
			"011011" when smallx = "0010011" and smally = "0001011" else
			"011011" when smallx = "0010100" and smally = "0001011" else
			"011011" when smallx = "0010101" and smally = "0001011" else
			"011011" when smallx = "0000000" and smally = "0001100" else
			"011011" when smallx = "0000001" and smally = "0001100" else
			"000000" when smallx = "0000010" and smally = "0001100" else
			"000000" when smallx = "0000011" and smally = "0001100" else
			"000000" when smallx = "0000100" and smally = "0001100" else
			"000000" when smallx = "0000101" and smally = "0001100" else
			"011011" when smallx = "0000110" and smally = "0001100" else
			"011011" when smallx = "0000111" and smally = "0001100" else
			"011011" when smallx = "0001000" and smally = "0001100" else
			"011011" when smallx = "0001001" and smally = "0001100" else
			"011011" when smallx = "0001010" and smally = "0001100" else
			"000000" when smallx = "0001011" and smally = "0001100" else
			"000000" when smallx = "0001100" and smally = "0001100" else
			"000000" when smallx = "0001101" and smally = "0001100" else
			"000000" when smallx = "0001110" and smally = "0001100" else
			"011011" when smallx = "0001111" and smally = "0001100" else
			"011011" when smallx = "0010000" and smally = "0001100" else
			"011011" when smallx = "0010001" and smally = "0001100" else
			"011011" when smallx = "0010010" and smally = "0001100" else
			"011011" when smallx = "0010011" and smally = "0001100" else
			"011011" when smallx = "0010100" and smally = "0001100" else
			"011011" when smallx = "0010101" and smally = "0001100" else
			"011011";
end if;
end process;
end;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity startscreen is
        port (
                x : in unsigned(9 downto 0); -- 5bit for 32 pixel bird
                y : in unsigned(9 downto 0);
                rgb : out std_logic_vector(5 downto 0);
				clk : in std_logic
        );
end startscreen;

architecture synth of startscreen is
        signal smallx : unsigned(6 downto 0);
        signal smally : unsigned(6 downto 0);
begin
        smallx <= x(9 downto 3); -- divide to get image size (16x16)
        smally <= y(9 downto 3);

process(clk) begin
if rising_edge(clk) then
        rgb <=
			"010000" when smallx = "0000100" and smally = "0000100" else
			"010000" when smallx = "0000101" and smally = "0000100" else
			"010000" when smallx = "0000110" and smally = "0000100" else
			"010000" when smallx = "0000111" and smally = "0000100" else
			"010000" when smallx = "0001000" and smally = "0000100" else
			"010000" when smallx = "0001001" and smally = "0000100" else
			"010000" when smallx = "0001010" and smally = "0000100" else
			"010000" when smallx = "0001011" and smally = "0000100" else
			"010000" when smallx = "0001100" and smally = "0000100" else
			"010000" when smallx = "0001101" and smally = "0000100" else
			"010000" when smallx = "0001110" and smally = "0000100" else
			"010000" when smallx = "0001111" and smally = "0000100" else
			"010000" when smallx = "0010000" and smally = "0000100" else
			"010000" when smallx = "0010001" and smally = "0000100" else
			"010000" when smallx = "0010010" and smally = "0000100" else
			"010000" when smallx = "0010011" and smally = "0000100" else
			"010000" when smallx = "0010100" and smally = "0000100" else
			"010000" when smallx = "0010101" and smally = "0000100" else
			"010000" when smallx = "0010110" and smally = "0000100" else
			"010000" when smallx = "0010111" and smally = "0000100" else
			"010000" when smallx = "0011000" and smally = "0000100" else
			"010000" when smallx = "0011001" and smally = "0000100" else
			"010000" when smallx = "0011010" and smally = "0000100" else
			"010000" when smallx = "0011011" and smally = "0000100" else
			"010000" when smallx = "0011100" and smally = "0000100" else
			"010000" when smallx = "0011101" and smally = "0000100" else
			"010000" when smallx = "0011110" and smally = "0000100" else
			"010000" when smallx = "0011111" and smally = "0000100" else
			"010000" when smallx = "0100000" and smally = "0000100" else
			"010000" when smallx = "0100001" and smally = "0000100" else
			"010000" when smallx = "0100010" and smally = "0000100" else
			"010000" when smallx = "0100011" and smally = "0000100" else
			"010000" when smallx = "0100100" and smally = "0000100" else
			"010000" when smallx = "0100101" and smally = "0000100" else
			"010000" when smallx = "0100110" and smally = "0000100" else
			"010000" when smallx = "0100111" and smally = "0000100" else
			"010000" when smallx = "0101000" and smally = "0000100" else
			"010000" when smallx = "0101001" and smally = "0000100" else
			"010000" when smallx = "0101010" and smally = "0000100" else
			"010000" when smallx = "0101011" and smally = "0000100" else
			"010000" when smallx = "0101100" and smally = "0000100" else
			"010000" when smallx = "0101101" and smally = "0000100" else
			"010000" when smallx = "0101110" and smally = "0000100" else
			"010000" when smallx = "0101111" and smally = "0000100" else
			"010000" when smallx = "0110000" and smally = "0000100" else
			"010000" when smallx = "0110001" and smally = "0000100" else
			"010000" when smallx = "0110010" and smally = "0000100" else
			"010000" when smallx = "0110011" and smally = "0000100" else
			"010000" when smallx = "0110100" and smally = "0000100" else
			"010000" when smallx = "0110101" and smally = "0000100" else
			"010000" when smallx = "0110110" and smally = "0000100" else
			"010000" when smallx = "0110111" and smally = "0000100" else
			"010000" when smallx = "0111000" and smally = "0000100" else
			"010000" when smallx = "0111001" and smally = "0000100" else
			"010000" when smallx = "0111010" and smally = "0000100" else
			"010000" when smallx = "0111011" and smally = "0000100" else
			"010000" when smallx = "0111100" and smally = "0000100" else
			"010000" when smallx = "0111101" and smally = "0000100" else
			"010000" when smallx = "0111110" and smally = "0000100" else
			"010000" when smallx = "0111111" and smally = "0000100" else
			"010000" when smallx = "1000000" and smally = "0000100" else
			"010000" when smallx = "1000001" and smally = "0000100" else
			"010000" when smallx = "1000010" and smally = "0000100" else
			"010000" when smallx = "1000011" and smally = "0000100" else
			"010000" when smallx = "1000100" and smally = "0000100" else
			"010000" when smallx = "1000101" and smally = "0000100" else
			"010000" when smallx = "1000110" and smally = "0000100" else
			"010000" when smallx = "1000111" and smally = "0000100" else
			"010000" when smallx = "1001000" and smally = "0000100" else
			"010000" when smallx = "1001001" and smally = "0000100" else
			"010000" when smallx = "1001010" and smally = "0000100" else
			"010000" when smallx = "0000100" and smally = "0000101" else
			"010000" when smallx = "0000101" and smally = "0000101" else
			"010000" when smallx = "0000110" and smally = "0000101" else
			"010000" when smallx = "0000111" and smally = "0000101" else
			"010000" when smallx = "0001000" and smally = "0000101" else
			"010000" when smallx = "0001001" and smally = "0000101" else
			"010000" when smallx = "0001010" and smally = "0000101" else
			"010000" when smallx = "0001011" and smally = "0000101" else
			"010000" when smallx = "0001100" and smally = "0000101" else
			"010000" when smallx = "0001101" and smally = "0000101" else
			"010000" when smallx = "0001110" and smally = "0000101" else
			"010000" when smallx = "0001111" and smally = "0000101" else
			"010000" when smallx = "0010000" and smally = "0000101" else
			"010000" when smallx = "0010001" and smally = "0000101" else
			"010000" when smallx = "0010010" and smally = "0000101" else
			"010000" when smallx = "0010011" and smally = "0000101" else
			"010000" when smallx = "0010100" and smally = "0000101" else
			"010000" when smallx = "0010101" and smally = "0000101" else
			"010000" when smallx = "0010110" and smally = "0000101" else
			"010000" when smallx = "0010111" and smally = "0000101" else
			"010000" when smallx = "0011000" and smally = "0000101" else
			"010000" when smallx = "0011001" and smally = "0000101" else
			"010000" when smallx = "0011010" and smally = "0000101" else
			"010000" when smallx = "0011011" and smally = "0000101" else
			"010000" when smallx = "0011100" and smally = "0000101" else
			"010000" when smallx = "0011101" and smally = "0000101" else
			"010000" when smallx = "0011110" and smally = "0000101" else
			"010000" when smallx = "0011111" and smally = "0000101" else
			"010000" when smallx = "0100000" and smally = "0000101" else
			"010000" when smallx = "0100001" and smally = "0000101" else
			"010000" when smallx = "0100010" and smally = "0000101" else
			"010000" when smallx = "0100011" and smally = "0000101" else
			"010000" when smallx = "0100100" and smally = "0000101" else
			"010000" when smallx = "0100101" and smally = "0000101" else
			"010000" when smallx = "0100110" and smally = "0000101" else
			"010000" when smallx = "0100111" and smally = "0000101" else
			"010000" when smallx = "0101000" and smally = "0000101" else
			"010000" when smallx = "0101001" and smally = "0000101" else
			"010000" when smallx = "0101010" and smally = "0000101" else
			"010000" when smallx = "0101011" and smally = "0000101" else
			"010000" when smallx = "0101100" and smally = "0000101" else
			"010000" when smallx = "0101101" and smally = "0000101" else
			"010000" when smallx = "0101110" and smally = "0000101" else
			"010000" when smallx = "0101111" and smally = "0000101" else
			"010000" when smallx = "0110000" and smally = "0000101" else
			"010000" when smallx = "0110001" and smally = "0000101" else
			"010000" when smallx = "0110010" and smally = "0000101" else
			"010000" when smallx = "0110011" and smally = "0000101" else
			"010000" when smallx = "0110100" and smally = "0000101" else
			"010000" when smallx = "0110101" and smally = "0000101" else
			"010000" when smallx = "0110110" and smally = "0000101" else
			"010000" when smallx = "0110111" and smally = "0000101" else
			"010000" when smallx = "0111000" and smally = "0000101" else
			"010000" when smallx = "0111001" and smally = "0000101" else
			"010000" when smallx = "0111010" and smally = "0000101" else
			"010000" when smallx = "0111011" and smally = "0000101" else
			"010000" when smallx = "0111100" and smally = "0000101" else
			"010000" when smallx = "0111101" and smally = "0000101" else
			"010000" when smallx = "0111110" and smally = "0000101" else
			"010000" when smallx = "0111111" and smally = "0000101" else
			"010000" when smallx = "1000000" and smally = "0000101" else
			"010000" when smallx = "1000001" and smally = "0000101" else
			"010000" when smallx = "1000010" and smally = "0000101" else
			"010000" when smallx = "1000011" and smally = "0000101" else
			"010000" when smallx = "1000100" and smally = "0000101" else
			"010000" when smallx = "1000101" and smally = "0000101" else
			"010000" when smallx = "1000110" and smally = "0000101" else
			"010000" when smallx = "1000111" and smally = "0000101" else
			"010000" when smallx = "1001000" and smally = "0000101" else
			"010000" when smallx = "1001001" and smally = "0000101" else
			"010000" when smallx = "1001010" and smally = "0000101" else
			"010000" when smallx = "0000100" and smally = "0000110" else
			"010000" when smallx = "0000101" and smally = "0000110" else
			"010000" when smallx = "0000110" and smally = "0000110" else
			"010000" when smallx = "0000111" and smally = "0000110" else
			"010000" when smallx = "0001000" and smally = "0000110" else
			"010000" when smallx = "0001001" and smally = "0000110" else
			"010000" when smallx = "0001010" and smally = "0000110" else
			"010000" when smallx = "0001011" and smally = "0000110" else
			"010000" when smallx = "0001100" and smally = "0000110" else
			"010000" when smallx = "0001101" and smally = "0000110" else
			"010000" when smallx = "0001110" and smally = "0000110" else
			"010000" when smallx = "0001111" and smally = "0000110" else
			"010000" when smallx = "0010000" and smally = "0000110" else
			"010000" when smallx = "0010001" and smally = "0000110" else
			"010000" when smallx = "0010010" and smally = "0000110" else
			"010000" when smallx = "0010011" and smally = "0000110" else
			"010000" when smallx = "0010100" and smally = "0000110" else
			"010000" when smallx = "0010101" and smally = "0000110" else
			"010000" when smallx = "0010110" and smally = "0000110" else
			"010000" when smallx = "0010111" and smally = "0000110" else
			"010000" when smallx = "0011000" and smally = "0000110" else
			"010000" when smallx = "0011001" and smally = "0000110" else
			"010000" when smallx = "0011010" and smally = "0000110" else
			"010000" when smallx = "0011011" and smally = "0000110" else
			"010000" when smallx = "0011100" and smally = "0000110" else
			"010000" when smallx = "0011101" and smally = "0000110" else
			"010000" when smallx = "0011110" and smally = "0000110" else
			"010000" when smallx = "0011111" and smally = "0000110" else
			"010000" when smallx = "0100000" and smally = "0000110" else
			"010000" when smallx = "0100001" and smally = "0000110" else
			"010000" when smallx = "0100010" and smally = "0000110" else
			"010000" when smallx = "0100011" and smally = "0000110" else
			"010000" when smallx = "0100100" and smally = "0000110" else
			"010000" when smallx = "0100101" and smally = "0000110" else
			"010000" when smallx = "0100110" and smally = "0000110" else
			"010000" when smallx = "0100111" and smally = "0000110" else
			"010000" when smallx = "0101000" and smally = "0000110" else
			"010000" when smallx = "0101001" and smally = "0000110" else
			"010000" when smallx = "0101010" and smally = "0000110" else
			"010000" when smallx = "0101011" and smally = "0000110" else
			"010000" when smallx = "0101100" and smally = "0000110" else
			"010000" when smallx = "0101101" and smally = "0000110" else
			"010000" when smallx = "0101110" and smally = "0000110" else
			"010000" when smallx = "0101111" and smally = "0000110" else
			"010000" when smallx = "0110000" and smally = "0000110" else
			"010000" when smallx = "0110001" and smally = "0000110" else
			"010000" when smallx = "0110010" and smally = "0000110" else
			"010000" when smallx = "0110011" and smally = "0000110" else
			"010000" when smallx = "0110100" and smally = "0000110" else
			"010000" when smallx = "0110101" and smally = "0000110" else
			"010000" when smallx = "0110110" and smally = "0000110" else
			"010000" when smallx = "0110111" and smally = "0000110" else
			"010000" when smallx = "0111000" and smally = "0000110" else
			"010000" when smallx = "0111001" and smally = "0000110" else
			"010000" when smallx = "0111010" and smally = "0000110" else
			"010000" when smallx = "0111011" and smally = "0000110" else
			"010000" when smallx = "0111100" and smally = "0000110" else
			"010000" when smallx = "0111101" and smally = "0000110" else
			"010000" when smallx = "0111110" and smally = "0000110" else
			"010000" when smallx = "0111111" and smally = "0000110" else
			"010000" when smallx = "1000000" and smally = "0000110" else
			"010000" when smallx = "1000001" and smally = "0000110" else
			"010000" when smallx = "1000010" and smally = "0000110" else
			"010000" when smallx = "1000011" and smally = "0000110" else
			"010000" when smallx = "1000100" and smally = "0000110" else
			"010000" when smallx = "1000101" and smally = "0000110" else
			"010000" when smallx = "1000110" and smally = "0000110" else
			"010000" when smallx = "1000111" and smally = "0000110" else
			"010000" when smallx = "1001000" and smally = "0000110" else
			"010000" when smallx = "1001001" and smally = "0000110" else
			"010000" when smallx = "1001010" and smally = "0000110" else
			"010000" when smallx = "0000100" and smally = "0000111" else
			"010000" when smallx = "0000101" and smally = "0000111" else
			"010000" when smallx = "0000110" and smally = "0000111" else
			"010000" when smallx = "0000111" and smally = "0000111" else
			"010000" when smallx = "0001000" and smally = "0000111" else
			"010000" when smallx = "0001001" and smally = "0000111" else
			"010000" when smallx = "0001010" and smally = "0000111" else
			"010000" when smallx = "0001011" and smally = "0000111" else
			"010000" when smallx = "0001100" and smally = "0000111" else
			"111111" when smallx = "0001101" and smally = "0000111" else
			"111111" when smallx = "0001110" and smally = "0000111" else
			"111111" when smallx = "0001111" and smally = "0000111" else
			"111111" when smallx = "0010000" and smally = "0000111" else
			"010000" when smallx = "0010001" and smally = "0000111" else
			"111111" when smallx = "0010010" and smally = "0000111" else
			"010000" when smallx = "0010011" and smally = "0000111" else
			"010000" when smallx = "0010100" and smally = "0000111" else
			"010000" when smallx = "0010101" and smally = "0000111" else
			"010000" when smallx = "0010110" and smally = "0000111" else
			"010000" when smallx = "0010111" and smally = "0000111" else
			"111111" when smallx = "0011000" and smally = "0000111" else
			"111111" when smallx = "0011001" and smally = "0000111" else
			"010000" when smallx = "0011010" and smally = "0000111" else
			"010000" when smallx = "0011011" and smally = "0000111" else
			"111111" when smallx = "0011100" and smally = "0000111" else
			"111111" when smallx = "0011101" and smally = "0000111" else
			"111111" when smallx = "0011110" and smally = "0000111" else
			"010000" when smallx = "0011111" and smally = "0000111" else
			"010000" when smallx = "0100000" and smally = "0000111" else
			"111111" when smallx = "0100001" and smally = "0000111" else
			"111111" when smallx = "0100010" and smally = "0000111" else
			"111111" when smallx = "0100011" and smally = "0000111" else
			"010000" when smallx = "0100100" and smally = "0000111" else
			"010000" when smallx = "0100101" and smally = "0000111" else
			"111111" when smallx = "0100110" and smally = "0000111" else
			"010000" when smallx = "0100111" and smally = "0000111" else
			"010000" when smallx = "0101000" and smally = "0000111" else
			"010000" when smallx = "0101001" and smally = "0000111" else
			"111111" when smallx = "0101010" and smally = "0000111" else
			"010000" when smallx = "0101011" and smally = "0000111" else
			"010000" when smallx = "0101100" and smally = "0000111" else
			"010000" when smallx = "0101101" and smally = "0000111" else
			"010000" when smallx = "0101110" and smally = "0000111" else
			"111111" when smallx = "0101111" and smally = "0000111" else
			"010000" when smallx = "0110000" and smally = "0000111" else
			"010000" when smallx = "0110001" and smally = "0000111" else
			"111111" when smallx = "0110010" and smally = "0000111" else
			"111111" when smallx = "0110011" and smally = "0000111" else
			"111111" when smallx = "0110100" and smally = "0000111" else
			"010000" when smallx = "0110101" and smally = "0000111" else
			"010000" when smallx = "0110110" and smally = "0000111" else
			"010000" when smallx = "0110111" and smally = "0000111" else
			"111111" when smallx = "0111000" and smally = "0000111" else
			"111111" when smallx = "0111001" and smally = "0000111" else
			"010000" when smallx = "0111010" and smally = "0000111" else
			"010000" when smallx = "0111011" and smally = "0000111" else
			"010000" when smallx = "0111100" and smally = "0000111" else
			"111111" when smallx = "0111101" and smally = "0000111" else
			"111111" when smallx = "0111110" and smally = "0000111" else
			"111111" when smallx = "0111111" and smally = "0000111" else
			"010000" when smallx = "1000000" and smally = "0000111" else
			"010000" when smallx = "1000001" and smally = "0000111" else
			"010000" when smallx = "1000010" and smally = "0000111" else
			"010000" when smallx = "1000011" and smally = "0000111" else
			"010000" when smallx = "1000100" and smally = "0000111" else
			"010000" when smallx = "1000101" and smally = "0000111" else
			"010000" when smallx = "1000110" and smally = "0000111" else
			"010000" when smallx = "1000111" and smally = "0000111" else
			"010000" when smallx = "1001000" and smally = "0000111" else
			"010000" when smallx = "1001001" and smally = "0000111" else
			"010000" when smallx = "1001010" and smally = "0000111" else
			"010000" when smallx = "0000100" and smally = "0001000" else
			"010000" when smallx = "0000101" and smally = "0001000" else
			"010000" when smallx = "0000110" and smally = "0001000" else
			"010000" when smallx = "0000111" and smally = "0001000" else
			"010000" when smallx = "0001000" and smally = "0001000" else
			"010000" when smallx = "0001001" and smally = "0001000" else
			"010000" when smallx = "0001010" and smally = "0001000" else
			"010000" when smallx = "0001011" and smally = "0001000" else
			"010000" when smallx = "0001100" and smally = "0001000" else
			"111111" when smallx = "0001101" and smally = "0001000" else
			"010000" when smallx = "0001110" and smally = "0001000" else
			"010000" when smallx = "0001111" and smally = "0001000" else
			"010000" when smallx = "0010000" and smally = "0001000" else
			"010000" when smallx = "0010001" and smally = "0001000" else
			"111111" when smallx = "0010010" and smally = "0001000" else
			"010000" when smallx = "0010011" and smally = "0001000" else
			"010000" when smallx = "0010100" and smally = "0001000" else
			"010000" when smallx = "0010101" and smally = "0001000" else
			"010000" when smallx = "0010110" and smally = "0001000" else
			"111111" when smallx = "0010111" and smally = "0001000" else
			"010000" when smallx = "0011000" and smally = "0001000" else
			"010000" when smallx = "0011001" and smally = "0001000" else
			"111111" when smallx = "0011010" and smally = "0001000" else
			"010000" when smallx = "0011011" and smally = "0001000" else
			"111111" when smallx = "0011100" and smally = "0001000" else
			"010000" when smallx = "0011101" and smally = "0001000" else
			"010000" when smallx = "0011110" and smally = "0001000" else
			"111111" when smallx = "0011111" and smally = "0001000" else
			"010000" when smallx = "0100000" and smally = "0001000" else
			"111111" when smallx = "0100001" and smally = "0001000" else
			"010000" when smallx = "0100010" and smally = "0001000" else
			"010000" when smallx = "0100011" and smally = "0001000" else
			"111111" when smallx = "0100100" and smally = "0001000" else
			"010000" when smallx = "0100101" and smally = "0001000" else
			"111111" when smallx = "0100110" and smally = "0001000" else
			"010000" when smallx = "0100111" and smally = "0001000" else
			"010000" when smallx = "0101000" and smally = "0001000" else
			"010000" when smallx = "0101001" and smally = "0001000" else
			"111111" when smallx = "0101010" and smally = "0001000" else
			"010000" when smallx = "0101011" and smally = "0001000" else
			"010000" when smallx = "0101100" and smally = "0001000" else
			"010000" when smallx = "0101101" and smally = "0001000" else
			"010000" when smallx = "0101110" and smally = "0001000" else
			"111111" when smallx = "0101111" and smally = "0001000" else
			"010000" when smallx = "0110000" and smally = "0001000" else
			"010000" when smallx = "0110001" and smally = "0001000" else
			"111111" when smallx = "0110010" and smally = "0001000" else
			"010000" when smallx = "0110011" and smally = "0001000" else
			"010000" when smallx = "0110100" and smally = "0001000" else
			"111111" when smallx = "0110101" and smally = "0001000" else
			"010000" when smallx = "0110110" and smally = "0001000" else
			"111111" when smallx = "0110111" and smally = "0001000" else
			"010000" when smallx = "0111000" and smally = "0001000" else
			"010000" when smallx = "0111001" and smally = "0001000" else
			"111111" when smallx = "0111010" and smally = "0001000" else
			"010000" when smallx = "0111011" and smally = "0001000" else
			"111111" when smallx = "0111100" and smally = "0001000" else
			"010000" when smallx = "0111101" and smally = "0001000" else
			"010000" when smallx = "0111110" and smally = "0001000" else
			"010000" when smallx = "0111111" and smally = "0001000" else
			"010000" when smallx = "1000000" and smally = "0001000" else
			"010000" when smallx = "1000001" and smally = "0001000" else
			"010000" when smallx = "1000010" and smally = "0001000" else
			"010000" when smallx = "1000011" and smally = "0001000" else
			"010000" when smallx = "1000100" and smally = "0001000" else
			"010000" when smallx = "1000101" and smally = "0001000" else
			"010000" when smallx = "1000110" and smally = "0001000" else
			"010000" when smallx = "1000111" and smally = "0001000" else
			"010000" when smallx = "1001000" and smally = "0001000" else
			"010000" when smallx = "1001001" and smally = "0001000" else
			"010000" when smallx = "1001010" and smally = "0001000" else
			"010000" when smallx = "0000100" and smally = "0001001" else
			"010000" when smallx = "0000101" and smally = "0001001" else
			"010000" when smallx = "0000110" and smally = "0001001" else
			"010000" when smallx = "0000111" and smally = "0001001" else
			"010000" when smallx = "0001000" and smally = "0001001" else
			"010000" when smallx = "0001001" and smally = "0001001" else
			"010000" when smallx = "0001010" and smally = "0001001" else
			"010000" when smallx = "0001011" and smally = "0001001" else
			"010000" when smallx = "0001100" and smally = "0001001" else
			"111111" when smallx = "0001101" and smally = "0001001" else
			"111111" when smallx = "0001110" and smally = "0001001" else
			"111111" when smallx = "0001111" and smally = "0001001" else
			"010000" when smallx = "0010000" and smally = "0001001" else
			"010000" when smallx = "0010001" and smally = "0001001" else
			"111111" when smallx = "0010010" and smally = "0001001" else
			"010000" when smallx = "0010011" and smally = "0001001" else
			"010000" when smallx = "0010100" and smally = "0001001" else
			"010000" when smallx = "0010101" and smally = "0001001" else
			"010000" when smallx = "0010110" and smally = "0001001" else
			"111111" when smallx = "0010111" and smally = "0001001" else
			"111111" when smallx = "0011000" and smally = "0001001" else
			"111111" when smallx = "0011001" and smally = "0001001" else
			"111111" when smallx = "0011010" and smally = "0001001" else
			"010000" when smallx = "0011011" and smally = "0001001" else
			"111111" when smallx = "0011100" and smally = "0001001" else
			"111111" when smallx = "0011101" and smally = "0001001" else
			"111111" when smallx = "0011110" and smally = "0001001" else
			"010000" when smallx = "0011111" and smally = "0001001" else
			"010000" when smallx = "0100000" and smally = "0001001" else
			"111111" when smallx = "0100001" and smally = "0001001" else
			"111111" when smallx = "0100010" and smally = "0001001" else
			"111111" when smallx = "0100011" and smally = "0001001" else
			"010000" when smallx = "0100100" and smally = "0001001" else
			"010000" when smallx = "0100101" and smally = "0001001" else
			"010000" when smallx = "0100110" and smally = "0001001" else
			"111111" when smallx = "0100111" and smally = "0001001" else
			"111111" when smallx = "0101000" and smally = "0001001" else
			"111111" when smallx = "0101001" and smally = "0001001" else
			"010000" when smallx = "0101010" and smally = "0001001" else
			"010000" when smallx = "0101011" and smally = "0001001" else
			"010000" when smallx = "0101100" and smally = "0001001" else
			"010000" when smallx = "0101101" and smally = "0001001" else
			"010000" when smallx = "0101110" and smally = "0001001" else
			"010000" when smallx = "0101111" and smally = "0001001" else
			"010000" when smallx = "0110000" and smally = "0001001" else
			"010000" when smallx = "0110001" and smally = "0001001" else
			"111111" when smallx = "0110010" and smally = "0001001" else
			"111111" when smallx = "0110011" and smally = "0001001" else
			"111111" when smallx = "0110100" and smally = "0001001" else
			"010000" when smallx = "0110101" and smally = "0001001" else
			"010000" when smallx = "0110110" and smally = "0001001" else
			"111111" when smallx = "0110111" and smally = "0001001" else
			"010000" when smallx = "0111000" and smally = "0001001" else
			"010000" when smallx = "0111001" and smally = "0001001" else
			"111111" when smallx = "0111010" and smally = "0001001" else
			"010000" when smallx = "0111011" and smally = "0001001" else
			"010000" when smallx = "0111100" and smally = "0001001" else
			"111111" when smallx = "0111101" and smally = "0001001" else
			"111111" when smallx = "0111110" and smally = "0001001" else
			"010000" when smallx = "0111111" and smally = "0001001" else
			"010000" when smallx = "1000000" and smally = "0001001" else
			"010000" when smallx = "1000001" and smally = "0001001" else
			"010000" when smallx = "1000010" and smally = "0001001" else
			"010000" when smallx = "1000011" and smally = "0001001" else
			"010000" when smallx = "1000100" and smally = "0001001" else
			"010000" when smallx = "1000101" and smally = "0001001" else
			"010000" when smallx = "1000110" and smally = "0001001" else
			"010000" when smallx = "1000111" and smally = "0001001" else
			"010000" when smallx = "1001000" and smally = "0001001" else
			"010000" when smallx = "1001001" and smally = "0001001" else
			"010000" when smallx = "1001010" and smally = "0001001" else
			"010000" when smallx = "0000100" and smally = "0001010" else
			"010000" when smallx = "0000101" and smally = "0001010" else
			"010000" when smallx = "0000110" and smally = "0001010" else
			"010000" when smallx = "0000111" and smally = "0001010" else
			"010000" when smallx = "0001000" and smally = "0001010" else
			"010000" when smallx = "0001001" and smally = "0001010" else
			"010000" when smallx = "0001010" and smally = "0001010" else
			"010000" when smallx = "0001011" and smally = "0001010" else
			"010000" when smallx = "0001100" and smally = "0001010" else
			"111111" when smallx = "0001101" and smally = "0001010" else
			"010000" when smallx = "0001110" and smally = "0001010" else
			"010000" when smallx = "0001111" and smally = "0001010" else
			"010000" when smallx = "0010000" and smally = "0001010" else
			"010000" when smallx = "0010001" and smally = "0001010" else
			"111111" when smallx = "0010010" and smally = "0001010" else
			"010000" when smallx = "0010011" and smally = "0001010" else
			"010000" when smallx = "0010100" and smally = "0001010" else
			"010000" when smallx = "0010101" and smally = "0001010" else
			"010000" when smallx = "0010110" and smally = "0001010" else
			"111111" when smallx = "0010111" and smally = "0001010" else
			"010000" when smallx = "0011000" and smally = "0001010" else
			"010000" when smallx = "0011001" and smally = "0001010" else
			"111111" when smallx = "0011010" and smally = "0001010" else
			"010000" when smallx = "0011011" and smally = "0001010" else
			"111111" when smallx = "0011100" and smally = "0001010" else
			"010000" when smallx = "0011101" and smally = "0001010" else
			"010000" when smallx = "0011110" and smally = "0001010" else
			"010000" when smallx = "0011111" and smally = "0001010" else
			"010000" when smallx = "0100000" and smally = "0001010" else
			"111111" when smallx = "0100001" and smally = "0001010" else
			"010000" when smallx = "0100010" and smally = "0001010" else
			"010000" when smallx = "0100011" and smally = "0001010" else
			"010000" when smallx = "0100100" and smally = "0001010" else
			"010000" when smallx = "0100101" and smally = "0001010" else
			"010000" when smallx = "0100110" and smally = "0001010" else
			"010000" when smallx = "0100111" and smally = "0001010" else
			"111111" when smallx = "0101000" and smally = "0001010" else
			"010000" when smallx = "0101001" and smally = "0001010" else
			"010000" when smallx = "0101010" and smally = "0001010" else
			"010000" when smallx = "0101011" and smally = "0001010" else
			"010000" when smallx = "0101100" and smally = "0001010" else
			"010000" when smallx = "0101101" and smally = "0001010" else
			"010000" when smallx = "0101110" and smally = "0001010" else
			"010000" when smallx = "0101111" and smally = "0001010" else
			"010000" when smallx = "0110000" and smally = "0001010" else
			"010000" when smallx = "0110001" and smally = "0001010" else
			"111111" when smallx = "0110010" and smally = "0001010" else
			"010000" when smallx = "0110011" and smally = "0001010" else
			"010000" when smallx = "0110100" and smally = "0001010" else
			"111111" when smallx = "0110101" and smally = "0001010" else
			"010000" when smallx = "0110110" and smally = "0001010" else
			"111111" when smallx = "0110111" and smally = "0001010" else
			"010000" when smallx = "0111000" and smally = "0001010" else
			"010000" when smallx = "0111001" and smally = "0001010" else
			"111111" when smallx = "0111010" and smally = "0001010" else
			"010000" when smallx = "0111011" and smally = "0001010" else
			"010000" when smallx = "0111100" and smally = "0001010" else
			"010000" when smallx = "0111101" and smally = "0001010" else
			"010000" when smallx = "0111110" and smally = "0001010" else
			"111111" when smallx = "0111111" and smally = "0001010" else
			"010000" when smallx = "1000000" and smally = "0001010" else
			"010000" when smallx = "1000001" and smally = "0001010" else
			"010000" when smallx = "1000010" and smally = "0001010" else
			"010000" when smallx = "1000011" and smally = "0001010" else
			"010000" when smallx = "1000100" and smally = "0001010" else
			"010000" when smallx = "1000101" and smally = "0001010" else
			"010000" when smallx = "1000110" and smally = "0001010" else
			"010000" when smallx = "1000111" and smally = "0001010" else
			"010000" when smallx = "1001000" and smally = "0001010" else
			"010000" when smallx = "1001001" and smally = "0001010" else
			"010000" when smallx = "1001010" and smally = "0001010" else
			"010000" when smallx = "0000100" and smally = "0001011" else
			"010000" when smallx = "0000101" and smally = "0001011" else
			"010000" when smallx = "0000110" and smally = "0001011" else
			"010000" when smallx = "0000111" and smally = "0001011" else
			"010000" when smallx = "0001000" and smally = "0001011" else
			"010000" when smallx = "0001001" and smally = "0001011" else
			"010000" when smallx = "0001010" and smally = "0001011" else
			"010000" when smallx = "0001011" and smally = "0001011" else
			"010000" when smallx = "0001100" and smally = "0001011" else
			"111111" when smallx = "0001101" and smally = "0001011" else
			"010000" when smallx = "0001110" and smally = "0001011" else
			"010000" when smallx = "0001111" and smally = "0001011" else
			"010000" when smallx = "0010000" and smally = "0001011" else
			"010000" when smallx = "0010001" and smally = "0001011" else
			"111111" when smallx = "0010010" and smally = "0001011" else
			"111111" when smallx = "0010011" and smally = "0001011" else
			"111111" when smallx = "0010100" and smally = "0001011" else
			"111111" when smallx = "0010101" and smally = "0001011" else
			"010000" when smallx = "0010110" and smally = "0001011" else
			"111111" when smallx = "0010111" and smally = "0001011" else
			"010000" when smallx = "0011000" and smally = "0001011" else
			"010000" when smallx = "0011001" and smally = "0001011" else
			"111111" when smallx = "0011010" and smally = "0001011" else
			"010000" when smallx = "0011011" and smally = "0001011" else
			"111111" when smallx = "0011100" and smally = "0001011" else
			"010000" when smallx = "0011101" and smally = "0001011" else
			"010000" when smallx = "0011110" and smally = "0001011" else
			"010000" when smallx = "0011111" and smally = "0001011" else
			"010000" when smallx = "0100000" and smally = "0001011" else
			"111111" when smallx = "0100001" and smally = "0001011" else
			"010000" when smallx = "0100010" and smally = "0001011" else
			"010000" when smallx = "0100011" and smally = "0001011" else
			"010000" when smallx = "0100100" and smally = "0001011" else
			"010000" when smallx = "0100101" and smally = "0001011" else
			"010000" when smallx = "0100110" and smally = "0001011" else
			"010000" when smallx = "0100111" and smally = "0001011" else
			"111111" when smallx = "0101000" and smally = "0001011" else
			"010000" when smallx = "0101001" and smally = "0001011" else
			"010000" when smallx = "0101010" and smally = "0001011" else
			"010000" when smallx = "0101011" and smally = "0001011" else
			"010000" when smallx = "0101100" and smally = "0001011" else
			"010000" when smallx = "0101101" and smally = "0001011" else
			"010000" when smallx = "0101110" and smally = "0001011" else
			"010000" when smallx = "0101111" and smally = "0001011" else
			"010000" when smallx = "0110000" and smally = "0001011" else
			"010000" when smallx = "0110001" and smally = "0001011" else
			"111111" when smallx = "0110010" and smally = "0001011" else
			"111111" when smallx = "0110011" and smally = "0001011" else
			"111111" when smallx = "0110100" and smally = "0001011" else
			"010000" when smallx = "0110101" and smally = "0001011" else
			"010000" when smallx = "0110110" and smally = "0001011" else
			"010000" when smallx = "0110111" and smally = "0001011" else
			"111111" when smallx = "0111000" and smally = "0001011" else
			"111111" when smallx = "0111001" and smally = "0001011" else
			"010000" when smallx = "0111010" and smally = "0001011" else
			"010000" when smallx = "0111011" and smally = "0001011" else
			"111111" when smallx = "0111100" and smally = "0001011" else
			"111111" when smallx = "0111101" and smally = "0001011" else
			"111111" when smallx = "0111110" and smally = "0001011" else
			"010000" when smallx = "0111111" and smally = "0001011" else
			"010000" when smallx = "1000000" and smally = "0001011" else
			"010000" when smallx = "1000001" and smally = "0001011" else
			"010000" when smallx = "1000010" and smally = "0001011" else
			"010000" when smallx = "1000011" and smally = "0001011" else
			"010000" when smallx = "1000100" and smally = "0001011" else
			"010000" when smallx = "1000101" and smally = "0001011" else
			"010000" when smallx = "1000110" and smally = "0001011" else
			"010000" when smallx = "1000111" and smally = "0001011" else
			"010000" when smallx = "1001000" and smally = "0001011" else
			"010000" when smallx = "1001001" and smally = "0001011" else
			"010000" when smallx = "1001010" and smally = "0001011" else
			"010000" when smallx = "0000100" and smally = "0001100" else
			"010000" when smallx = "0000101" and smally = "0001100" else
			"010000" when smallx = "0000110" and smally = "0001100" else
			"010000" when smallx = "0000111" and smally = "0001100" else
			"010000" when smallx = "0001000" and smally = "0001100" else
			"010000" when smallx = "0001001" and smally = "0001100" else
			"010000" when smallx = "0001010" and smally = "0001100" else
			"010000" when smallx = "0001011" and smally = "0001100" else
			"010000" when smallx = "0001100" and smally = "0001100" else
			"010000" when smallx = "0001101" and smally = "0001100" else
			"010000" when smallx = "0001110" and smally = "0001100" else
			"010000" when smallx = "0001111" and smally = "0001100" else
			"010000" when smallx = "0010000" and smally = "0001100" else
			"010000" when smallx = "0010001" and smally = "0001100" else
			"010000" when smallx = "0010010" and smally = "0001100" else
			"010000" when smallx = "0010011" and smally = "0001100" else
			"010000" when smallx = "0010100" and smally = "0001100" else
			"010000" when smallx = "0010101" and smally = "0001100" else
			"010000" when smallx = "0010110" and smally = "0001100" else
			"010000" when smallx = "0010111" and smally = "0001100" else
			"010000" when smallx = "0011000" and smally = "0001100" else
			"010000" when smallx = "0011001" and smally = "0001100" else
			"010000" when smallx = "0011010" and smally = "0001100" else
			"010000" when smallx = "0011011" and smally = "0001100" else
			"010000" when smallx = "0011100" and smally = "0001100" else
			"010000" when smallx = "0011101" and smally = "0001100" else
			"010000" when smallx = "0011110" and smally = "0001100" else
			"010000" when smallx = "0011111" and smally = "0001100" else
			"010000" when smallx = "0100000" and smally = "0001100" else
			"010000" when smallx = "0100001" and smally = "0001100" else
			"010000" when smallx = "0100010" and smally = "0001100" else
			"010000" when smallx = "0100011" and smally = "0001100" else
			"010000" when smallx = "0100100" and smally = "0001100" else
			"010000" when smallx = "0100101" and smally = "0001100" else
			"010000" when smallx = "0100110" and smally = "0001100" else
			"010000" when smallx = "0100111" and smally = "0001100" else
			"010000" when smallx = "0101000" and smally = "0001100" else
			"010000" when smallx = "0101001" and smally = "0001100" else
			"010000" when smallx = "0101010" and smally = "0001100" else
			"010000" when smallx = "0101011" and smally = "0001100" else
			"010000" when smallx = "0101100" and smally = "0001100" else
			"010000" when smallx = "0101101" and smally = "0001100" else
			"010000" when smallx = "0101110" and smally = "0001100" else
			"010000" when smallx = "0101111" and smally = "0001100" else
			"010000" when smallx = "0110000" and smally = "0001100" else
			"010000" when smallx = "0110001" and smally = "0001100" else
			"010000" when smallx = "0110010" and smally = "0001100" else
			"010000" when smallx = "0110011" and smally = "0001100" else
			"010000" when smallx = "0110100" and smally = "0001100" else
			"010000" when smallx = "0110101" and smally = "0001100" else
			"010000" when smallx = "0110110" and smally = "0001100" else
			"010000" when smallx = "0110111" and smally = "0001100" else
			"010000" when smallx = "0111000" and smally = "0001100" else
			"010000" when smallx = "0111001" and smally = "0001100" else
			"010000" when smallx = "0111010" and smally = "0001100" else
			"010000" when smallx = "0111011" and smally = "0001100" else
			"010000" when smallx = "0111100" and smally = "0001100" else
			"010000" when smallx = "0111101" and smally = "0001100" else
			"010000" when smallx = "0111110" and smally = "0001100" else
			"010000" when smallx = "0111111" and smally = "0001100" else
			"010000" when smallx = "1000000" and smally = "0001100" else
			"010000" when smallx = "1000001" and smally = "0001100" else
			"010000" when smallx = "1000010" and smally = "0001100" else
			"010000" when smallx = "1000011" and smally = "0001100" else
			"010000" when smallx = "1000100" and smally = "0001100" else
			"010000" when smallx = "1000101" and smally = "0001100" else
			"010000" when smallx = "1000110" and smally = "0001100" else
			"010000" when smallx = "1000111" and smally = "0001100" else
			"010000" when smallx = "1001000" and smally = "0001100" else
			"010000" when smallx = "1001001" and smally = "0001100" else
			"010000" when smallx = "1001010" and smally = "0001100" else
			"010000" when smallx = "0000100" and smally = "0001101" else
			"010000" when smallx = "0000101" and smally = "0001101" else
			"010000" when smallx = "0000110" and smally = "0001101" else
			"010000" when smallx = "0000111" and smally = "0001101" else
			"010000" when smallx = "0001000" and smally = "0001101" else
			"010000" when smallx = "0001001" and smally = "0001101" else
			"010000" when smallx = "0001010" and smally = "0001101" else
			"010000" when smallx = "0001011" and smally = "0001101" else
			"010000" when smallx = "0001100" and smally = "0001101" else
			"010000" when smallx = "0001101" and smally = "0001101" else
			"010000" when smallx = "0001110" and smally = "0001101" else
			"010000" when smallx = "0001111" and smally = "0001101" else
			"010000" when smallx = "0010000" and smally = "0001101" else
			"010000" when smallx = "0010001" and smally = "0001101" else
			"010000" when smallx = "0010010" and smally = "0001101" else
			"010000" when smallx = "0010011" and smally = "0001101" else
			"010000" when smallx = "0010100" and smally = "0001101" else
			"010000" when smallx = "0010101" and smally = "0001101" else
			"010000" when smallx = "0010110" and smally = "0001101" else
			"010000" when smallx = "0010111" and smally = "0001101" else
			"010000" when smallx = "0011000" and smally = "0001101" else
			"010000" when smallx = "0011001" and smally = "0001101" else
			"010000" when smallx = "0011010" and smally = "0001101" else
			"010000" when smallx = "0011011" and smally = "0001101" else
			"010000" when smallx = "0011100" and smally = "0001101" else
			"010000" when smallx = "0011101" and smally = "0001101" else
			"010000" when smallx = "0011110" and smally = "0001101" else
			"010000" when smallx = "0011111" and smally = "0001101" else
			"010000" when smallx = "0100000" and smally = "0001101" else
			"010000" when smallx = "0100001" and smally = "0001101" else
			"010000" when smallx = "0100010" and smally = "0001101" else
			"010000" when smallx = "0100011" and smally = "0001101" else
			"010000" when smallx = "0100100" and smally = "0001101" else
			"010000" when smallx = "0100101" and smally = "0001101" else
			"010000" when smallx = "0100110" and smally = "0001101" else
			"010000" when smallx = "0100111" and smally = "0001101" else
			"010000" when smallx = "0101000" and smally = "0001101" else
			"010000" when smallx = "0101001" and smally = "0001101" else
			"010000" when smallx = "0101010" and smally = "0001101" else
			"010000" when smallx = "0101011" and smally = "0001101" else
			"010000" when smallx = "0101100" and smally = "0001101" else
			"010000" when smallx = "0101101" and smally = "0001101" else
			"010000" when smallx = "0101110" and smally = "0001101" else
			"010000" when smallx = "0101111" and smally = "0001101" else
			"010000" when smallx = "0110000" and smally = "0001101" else
			"010000" when smallx = "0110001" and smally = "0001101" else
			"010000" when smallx = "0110010" and smally = "0001101" else
			"010000" when smallx = "0110011" and smally = "0001101" else
			"010000" when smallx = "0110100" and smally = "0001101" else
			"010000" when smallx = "0110101" and smally = "0001101" else
			"010000" when smallx = "0110110" and smally = "0001101" else
			"010000" when smallx = "0110111" and smally = "0001101" else
			"010000" when smallx = "0111000" and smally = "0001101" else
			"010000" when smallx = "0111001" and smally = "0001101" else
			"010000" when smallx = "0111010" and smally = "0001101" else
			"010000" when smallx = "0111011" and smally = "0001101" else
			"010000" when smallx = "0111100" and smally = "0001101" else
			"010000" when smallx = "0111101" and smally = "0001101" else
			"010000" when smallx = "0111110" and smally = "0001101" else
			"010000" when smallx = "0111111" and smally = "0001101" else
			"010000" when smallx = "1000000" and smally = "0001101" else
			"010000" when smallx = "1000001" and smally = "0001101" else
			"010000" when smallx = "1000010" and smally = "0001101" else
			"010000" when smallx = "1000011" and smally = "0001101" else
			"010000" when smallx = "1000100" and smally = "0001101" else
			"010000" when smallx = "1000101" and smally = "0001101" else
			"010000" when smallx = "1000110" and smally = "0001101" else
			"010000" when smallx = "1000111" and smally = "0001101" else
			"010000" when smallx = "1001000" and smally = "0001101" else
			"010000" when smallx = "1001001" and smally = "0001101" else
			"010000" when smallx = "1001010" and smally = "0001101" else
			"010000" when smallx = "0000100" and smally = "0001110" else
			"010000" when smallx = "0000101" and smally = "0001110" else
			"010000" when smallx = "0000110" and smally = "0001110" else
			"010000" when smallx = "0000111" and smally = "0001110" else
			"010000" when smallx = "0001000" and smally = "0001110" else
			"010000" when smallx = "0001001" and smally = "0001110" else
			"010000" when smallx = "0001010" and smally = "0001110" else
			"010000" when smallx = "0001011" and smally = "0001110" else
			"010000" when smallx = "0001100" and smally = "0001110" else
			"010000" when smallx = "0001101" and smally = "0001110" else
			"010000" when smallx = "0001110" and smally = "0001110" else
			"010000" when smallx = "0001111" and smally = "0001110" else
			"010000" when smallx = "0010000" and smally = "0001110" else
			"010000" when smallx = "0010001" and smally = "0001110" else
			"010000" when smallx = "0010010" and smally = "0001110" else
			"010000" when smallx = "0010011" and smally = "0001110" else
			"010000" when smallx = "0010100" and smally = "0001110" else
			"010000" when smallx = "0010101" and smally = "0001110" else
			"010000" when smallx = "0010110" and smally = "0001110" else
			"010000" when smallx = "0010111" and smally = "0001110" else
			"010000" when smallx = "0011000" and smally = "0001110" else
			"010000" when smallx = "0011001" and smally = "0001110" else
			"010000" when smallx = "0011010" and smally = "0001110" else
			"010000" when smallx = "0011011" and smally = "0001110" else
			"010000" when smallx = "0011100" and smally = "0001110" else
			"010000" when smallx = "0011101" and smally = "0001110" else
			"010000" when smallx = "0011110" and smally = "0001110" else
			"010000" when smallx = "0011111" and smally = "0001110" else
			"010000" when smallx = "0100000" and smally = "0001110" else
			"010000" when smallx = "0100001" and smally = "0001110" else
			"010000" when smallx = "0100010" and smally = "0001110" else
			"010000" when smallx = "0100011" and smally = "0001110" else
			"010000" when smallx = "0100100" and smally = "0001110" else
			"010000" when smallx = "0100101" and smally = "0001110" else
			"010000" when smallx = "0100110" and smally = "0001110" else
			"010000" when smallx = "0100111" and smally = "0001110" else
			"010000" when smallx = "0101000" and smally = "0001110" else
			"010000" when smallx = "0101001" and smally = "0001110" else
			"010000" when smallx = "0101010" and smally = "0001110" else
			"010000" when smallx = "0101011" and smally = "0001110" else
			"010000" when smallx = "0101100" and smally = "0001110" else
			"010000" when smallx = "0101101" and smally = "0001110" else
			"010000" when smallx = "0101110" and smally = "0001110" else
			"010000" when smallx = "0101111" and smally = "0001110" else
			"010000" when smallx = "0110000" and smally = "0001110" else
			"010000" when smallx = "0110001" and smally = "0001110" else
			"010000" when smallx = "0110010" and smally = "0001110" else
			"010000" when smallx = "0110011" and smally = "0001110" else
			"010000" when smallx = "0110100" and smally = "0001110" else
			"010000" when smallx = "0110101" and smally = "0001110" else
			"010000" when smallx = "0110110" and smally = "0001110" else
			"010000" when smallx = "0110111" and smally = "0001110" else
			"010000" when smallx = "0111000" and smally = "0001110" else
			"010000" when smallx = "0111001" and smally = "0001110" else
			"010000" when smallx = "0111010" and smally = "0001110" else
			"010000" when smallx = "0111011" and smally = "0001110" else
			"010000" when smallx = "0111100" and smally = "0001110" else
			"010000" when smallx = "0111101" and smally = "0001110" else
			"010000" when smallx = "0111110" and smally = "0001110" else
			"010000" when smallx = "0111111" and smally = "0001110" else
			"010000" when smallx = "1000000" and smally = "0001110" else
			"010000" when smallx = "1000001" and smally = "0001110" else
			"010000" when smallx = "1000010" and smally = "0001110" else
			"010000" when smallx = "1000011" and smally = "0001110" else
			"010000" when smallx = "1000100" and smally = "0001110" else
			"010000" when smallx = "1000101" and smally = "0001110" else
			"010000" when smallx = "1000110" and smally = "0001110" else
			"010000" when smallx = "1000111" and smally = "0001110" else
			"010000" when smallx = "1001000" and smally = "0001110" else
			"010000" when smallx = "1001001" and smally = "0001110" else
			"010000" when smallx = "1001010" and smally = "0001110" else
			"111111" when smallx = "0010101" and smally = "0010011" else
			"111111" when smallx = "0010110" and smally = "0010011" else
			"111111" when smallx = "0010111" and smally = "0010011" else
			"111111" when smallx = "0011010" and smally = "0010011" else
			"111111" when smallx = "0011011" and smally = "0010011" else
			"111111" when smallx = "0011111" and smally = "0010011" else
			"111111" when smallx = "0100000" and smally = "0010011" else
			"111111" when smallx = "0100011" and smally = "0010011" else
			"111111" when smallx = "0100100" and smally = "0010011" else
			"111111" when smallx = "0100101" and smally = "0010011" else
			"111111" when smallx = "0101000" and smally = "0010011" else
			"111111" when smallx = "0101001" and smally = "0010011" else
			"111111" when smallx = "0101010" and smally = "0010011" else
			"111111" when smallx = "0101011" and smally = "0010011" else
			"111111" when smallx = "0010100" and smally = "0010100" else
			"111111" when smallx = "0011001" and smally = "0010100" else
			"111111" when smallx = "0011100" and smally = "0010100" else
			"111111" when smallx = "0011110" and smally = "0010100" else
			"111111" when smallx = "0100001" and smally = "0010100" else
			"111111" when smallx = "0100011" and smally = "0010100" else
			"111111" when smallx = "0100110" and smally = "0010100" else
			"111111" when smallx = "0101000" and smally = "0010100" else
			"111111" when smallx = "0101110" and smally = "0010100" else
			"111111" when smallx = "0010101" and smally = "0010101" else
			"111111" when smallx = "0010110" and smally = "0010101" else
			"111111" when smallx = "0011001" and smally = "0010101" else
			"111111" when smallx = "0011110" and smally = "0010101" else
			"111111" when smallx = "0100001" and smally = "0010101" else
			"111111" when smallx = "0100011" and smally = "0010101" else
			"111111" when smallx = "0100100" and smally = "0010101" else
			"111111" when smallx = "0100101" and smally = "0010101" else
			"111111" when smallx = "0101000" and smally = "0010101" else
			"111111" when smallx = "0101001" and smally = "0010101" else
			"111111" when smallx = "0101010" and smally = "0010101" else
			"111111" when smallx = "0010111" and smally = "0010110" else
			"111111" when smallx = "0011001" and smally = "0010110" else
			"111111" when smallx = "0011100" and smally = "0010110" else
			"111111" when smallx = "0011110" and smally = "0010110" else
			"111111" when smallx = "0100001" and smally = "0010110" else
			"111111" when smallx = "0100011" and smally = "0010110" else
			"111111" when smallx = "0100101" and smally = "0010110" else
			"111111" when smallx = "0101000" and smally = "0010110" else
			"111111" when smallx = "0101110" and smally = "0010110" else
			"111111" when smallx = "0010100" and smally = "0010111" else
			"111111" when smallx = "0010101" and smally = "0010111" else
			"111111" when smallx = "0010110" and smally = "0010111" else
			"111111" when smallx = "0011010" and smally = "0010111" else
			"111111" when smallx = "0011011" and smally = "0010111" else
			"111111" when smallx = "0011111" and smally = "0010111" else
			"111111" when smallx = "0100000" and smally = "0010111" else
			"111111" when smallx = "0100011" and smally = "0010111" else
			"111111" when smallx = "0100110" and smally = "0010111" else
			"111111" when smallx = "0101000" and smally = "0010111" else
			"111111" when smallx = "0101001" and smally = "0010111" else
			"111111" when smallx = "0101010" and smally = "0010111" else
			"111111" when smallx = "0101011" and smally = "0010111" else
			"000000" when smallx = "0100101" and smally = "0011110" else
			"000000" when smallx = "0100110" and smally = "0011110" else
			"000000" when smallx = "0100111" and smally = "0011110" else
			"000000" when smallx = "0101000" and smally = "0011110" else
			"000000" when smallx = "0101001" and smally = "0011110" else
			"000000" when smallx = "0101010" and smally = "0011110" else
			"000000" when smallx = "0101011" and smally = "0011110" else
			"000000" when smallx = "0101100" and smally = "0011110" else
			"000000" when smallx = "0100100" and smally = "0011111" else
			"010101" when smallx = "0100101" and smally = "0011111" else
			"010101" when smallx = "0100110" and smally = "0011111" else
			"010101" when smallx = "0100111" and smally = "0011111" else
			"010101" when smallx = "0101000" and smally = "0011111" else
			"010101" when smallx = "0101001" and smally = "0011111" else
			"000000" when smallx = "0101010" and smally = "0011111" else
			"101010" when smallx = "0101011" and smally = "0011111" else
			"101010" when smallx = "0101100" and smally = "0011111" else
			"000000" when smallx = "0101101" and smally = "0011111" else
			"000000" when smallx = "0100001" and smally = "0100000" else
			"000000" when smallx = "0100010" and smally = "0100000" else
			"000000" when smallx = "0100011" and smally = "0100000" else
			"000000" when smallx = "0100100" and smally = "0100000" else
			"010101" when smallx = "0100101" and smally = "0100000" else
			"010101" when smallx = "0100110" and smally = "0100000" else
			"010101" when smallx = "0100111" and smally = "0100000" else
			"010101" when smallx = "0101000" and smally = "0100000" else
			"010101" when smallx = "0101001" and smally = "0100000" else
			"000000" when smallx = "0101010" and smally = "0100000" else
			"101010" when smallx = "0101011" and smally = "0100000" else
			"101010" when smallx = "0101100" and smally = "0100000" else
			"101010" when smallx = "0101101" and smally = "0100000" else
			"000000" when smallx = "0101110" and smally = "0100000" else
			"000000" when smallx = "0100000" and smally = "0100001" else
			"101010" when smallx = "0100001" and smally = "0100001" else
			"101010" when smallx = "0100010" and smally = "0100001" else
			"101010" when smallx = "0100011" and smally = "0100001" else
			"101010" when smallx = "0100100" and smally = "0100001" else
			"000000" when smallx = "0100101" and smally = "0100001" else
			"010101" when smallx = "0100110" and smally = "0100001" else
			"010101" when smallx = "0100111" and smally = "0100001" else
			"010101" when smallx = "0101000" and smally = "0100001" else
			"000000" when smallx = "0101001" and smally = "0100001" else
			"101010" when smallx = "0101010" and smally = "0100001" else
			"101010" when smallx = "0101011" and smally = "0100001" else
			"101010" when smallx = "0101100" and smally = "0100001" else
			"101010" when smallx = "0101101" and smally = "0100001" else
			"000000" when smallx = "0101110" and smally = "0100001" else
			"000000" when smallx = "0011111" and smally = "0100010" else
			"101010" when smallx = "0100000" and smally = "0100010" else
			"101010" when smallx = "0100001" and smally = "0100010" else
			"101010" when smallx = "0100010" and smally = "0100010" else
			"101010" when smallx = "0100011" and smally = "0100010" else
			"101010" when smallx = "0100100" and smally = "0100010" else
			"101010" when smallx = "0100101" and smally = "0100010" else
			"000000" when smallx = "0100110" and smally = "0100010" else
			"000000" when smallx = "0100111" and smally = "0100010" else
			"000000" when smallx = "0101000" and smally = "0100010" else
			"101010" when smallx = "0101001" and smally = "0100010" else
			"101010" when smallx = "0101010" and smally = "0100010" else
			"101010" when smallx = "0101011" and smally = "0100010" else
			"101010" when smallx = "0101100" and smally = "0100010" else
			"101010" when smallx = "0101101" and smally = "0100010" else
			"000000" when smallx = "0101110" and smally = "0100010" else
			"000000" when smallx = "0011111" and smally = "0100011" else
			"101010" when smallx = "0100000" and smally = "0100011" else
			"101010" when smallx = "0100001" and smally = "0100011" else
			"101010" when smallx = "0100010" and smally = "0100011" else
			"101010" when smallx = "0100011" and smally = "0100011" else
			"101010" when smallx = "0100100" and smally = "0100011" else
			"101010" when smallx = "0100101" and smally = "0100011" else
			"101010" when smallx = "0100110" and smally = "0100011" else
			"101010" when smallx = "0100111" and smally = "0100011" else
			"101010" when smallx = "0101000" and smally = "0100011" else
			"101010" when smallx = "0101001" and smally = "0100011" else
			"101010" when smallx = "0101010" and smally = "0100011" else
			"101010" when smallx = "0101011" and smally = "0100011" else
			"000000" when smallx = "0101100" and smally = "0100011" else
			"101010" when smallx = "0101101" and smally = "0100011" else
			"000000" when smallx = "0101110" and smally = "0100011" else
			"000000" when smallx = "0110000" and smally = "0100011" else
			"000000" when smallx = "0110001" and smally = "0100011" else
			"000000" when smallx = "0011101" and smally = "0100100" else
			"000000" when smallx = "0011110" and smally = "0100100" else
			"000000" when smallx = "0011111" and smally = "0100100" else
			"101010" when smallx = "0100000" and smally = "0100100" else
			"101010" when smallx = "0100001" and smally = "0100100" else
			"101010" when smallx = "0100010" and smally = "0100100" else
			"101010" when smallx = "0100011" and smally = "0100100" else
			"101010" when smallx = "0100100" and smally = "0100100" else
			"101010" when smallx = "0100101" and smally = "0100100" else
			"101010" when smallx = "0100110" and smally = "0100100" else
			"101010" when smallx = "0100111" and smally = "0100100" else
			"101010" when smallx = "0101000" and smally = "0100100" else
			"101010" when smallx = "0101001" and smally = "0100100" else
			"101010" when smallx = "0101010" and smally = "0100100" else
			"101010" when smallx = "0101011" and smally = "0100100" else
			"101010" when smallx = "0101100" and smally = "0100100" else
			"101010" when smallx = "0101101" and smally = "0100100" else
			"000000" when smallx = "0101110" and smally = "0100100" else
			"000000" when smallx = "0101111" and smally = "0100100" else
			"101010" when smallx = "0110000" and smally = "0100100" else
			"101010" when smallx = "0110001" and smally = "0100100" else
			"000000" when smallx = "0110010" and smally = "0100100" else
			"000000" when smallx = "0011111" and smally = "0100101" else
			"101010" when smallx = "0100000" and smally = "0100101" else
			"101010" when smallx = "0100001" and smally = "0100101" else
			"101010" when smallx = "0100010" and smally = "0100101" else
			"101010" when smallx = "0100011" and smally = "0100101" else
			"101010" when smallx = "0100100" and smally = "0100101" else
			"101010" when smallx = "0100101" and smally = "0100101" else
			"101010" when smallx = "0100110" and smally = "0100101" else
			"101010" when smallx = "0100111" and smally = "0100101" else
			"101010" when smallx = "0101000" and smally = "0100101" else
			"101010" when smallx = "0101001" and smally = "0100101" else
			"101010" when smallx = "0101010" and smally = "0100101" else
			"101010" when smallx = "0101011" and smally = "0100101" else
			"101010" when smallx = "0101100" and smally = "0100101" else
			"101010" when smallx = "0101101" and smally = "0100101" else
			"101010" when smallx = "0101110" and smally = "0100101" else
			"101010" when smallx = "0101111" and smally = "0100101" else
			"101010" when smallx = "0110000" and smally = "0100101" else
			"000000" when smallx = "0110001" and smally = "0100101" else
			"000000" when smallx = "0011111" and smally = "0100110" else
			"101010" when smallx = "0100000" and smally = "0100110" else
			"101010" when smallx = "0100001" and smally = "0100110" else
			"000000" when smallx = "0100010" and smally = "0100110" else
			"000000" when smallx = "0100011" and smally = "0100110" else
			"000000" when smallx = "0100100" and smally = "0100110" else
			"000000" when smallx = "0100101" and smally = "0100110" else
			"000000" when smallx = "0100110" and smally = "0100110" else
			"000000" when smallx = "0100111" and smally = "0100110" else
			"000000" when smallx = "0101000" and smally = "0100110" else
			"101010" when smallx = "0101001" and smally = "0100110" else
			"101010" when smallx = "0101010" and smally = "0100110" else
			"101010" when smallx = "0101011" and smally = "0100110" else
			"101010" when smallx = "0101100" and smally = "0100110" else
			"101010" when smallx = "0101101" and smally = "0100110" else
			"000000" when smallx = "0101110" and smally = "0100110" else
			"000000" when smallx = "0101111" and smally = "0100110" else
			"000000" when smallx = "0110000" and smally = "0100110" else
			"000000" when smallx = "0011111" and smally = "0100111" else
			"101010" when smallx = "0100000" and smally = "0100111" else
			"101010" when smallx = "0100001" and smally = "0100111" else
			"000000" when smallx = "0100010" and smally = "0100111" else
			"000000" when smallx = "0101000" and smally = "0100111" else
			"101010" when smallx = "0101001" and smally = "0100111" else
			"101010" when smallx = "0101010" and smally = "0100111" else
			"000000" when smallx = "0101011" and smally = "0100111" else
			"000000" when smallx = "0101100" and smally = "0100111" else
			"000000" when smallx = "0101101" and smally = "0100111" else
			"000000" when smallx = "0011111" and smally = "0101000" else
			"101010" when smallx = "0100000" and smally = "0101000" else
			"101010" when smallx = "0100001" and smally = "0101000" else
			"000000" when smallx = "0100010" and smally = "0101000" else
			"000000" when smallx = "0101000" and smally = "0101000" else
			"101010" when smallx = "0101001" and smally = "0101000" else
			"101010" when smallx = "0101010" and smally = "0101000" else
			"000000" when smallx = "0101011" and smally = "0101000" else
			"000000" when smallx = "0011111" and smally = "0101001" else
			"101010" when smallx = "0100000" and smally = "0101001" else
			"101010" when smallx = "0100001" and smally = "0101001" else
			"000000" when smallx = "0100010" and smally = "0101001" else
			"000000" when smallx = "0101000" and smally = "0101001" else
			"101010" when smallx = "0101001" and smally = "0101001" else
			"101010" when smallx = "0101010" and smally = "0101001" else
			"000000" when smallx = "0101011" and smally = "0101001" else
			"000000" when smallx = "0011111" and smally = "0101010" else
			"000000" when smallx = "0100000" and smally = "0101010" else
			"000000" when smallx = "0100001" and smally = "0101010" else
			"000000" when smallx = "0100010" and smally = "0101010" else
			"000000" when smallx = "0101000" and smally = "0101010" else
			"000000" when smallx = "0101001" and smally = "0101010" else
			"000000" when smallx = "0101010" and smally = "0101010" else
			"000000" when smallx = "0101011" and smally = "0101010" else
			"111111" when smallx = "0001101" and smally = "0110010" else
			"111111" when smallx = "0001110" and smally = "0110010" else
			"111111" when smallx = "0001111" and smally = "0110010" else
			"111111" when smallx = "0010010" and smally = "0110010" else
			"111111" when smallx = "0010011" and smally = "0110010" else
			"111111" when smallx = "0010100" and smally = "0110010" else
			"111111" when smallx = "0010111" and smally = "0110010" else
			"111111" when smallx = "0011000" and smally = "0110010" else
			"111111" when smallx = "0011001" and smally = "0110010" else
			"111111" when smallx = "0011010" and smally = "0110010" else
			"111111" when smallx = "0011101" and smally = "0110010" else
			"111111" when smallx = "0011110" and smally = "0110010" else
			"111111" when smallx = "0011111" and smally = "0110010" else
			"111111" when smallx = "0100010" and smally = "0110010" else
			"111111" when smallx = "0100011" and smally = "0110010" else
			"111111" when smallx = "0100100" and smally = "0110010" else
			"111111" when smallx = "0101001" and smally = "0110010" else
			"111111" when smallx = "0101010" and smally = "0110010" else
			"111111" when smallx = "0101011" and smally = "0110010" else
			"111111" when smallx = "0101101" and smally = "0110010" else
			"111111" when smallx = "0101110" and smally = "0110010" else
			"111111" when smallx = "0101111" and smally = "0110010" else
			"111111" when smallx = "0110000" and smally = "0110010" else
			"111111" when smallx = "0110001" and smally = "0110010" else
			"111111" when smallx = "0110100" and smally = "0110010" else
			"111111" when smallx = "0110101" and smally = "0110010" else
			"111111" when smallx = "0111000" and smally = "0110010" else
			"111111" when smallx = "0111001" and smally = "0110010" else
			"111111" when smallx = "0111010" and smally = "0110010" else
			"111111" when smallx = "0111101" and smally = "0110010" else
			"111111" when smallx = "0111110" and smally = "0110010" else
			"111111" when smallx = "0111111" and smally = "0110010" else
			"111111" when smallx = "1000000" and smally = "0110010" else
			"111111" when smallx = "1000001" and smally = "0110010" else
			"111111" when smallx = "0001101" and smally = "0110011" else
			"111111" when smallx = "0010000" and smally = "0110011" else
			"111111" when smallx = "0010010" and smally = "0110011" else
			"111111" when smallx = "0010101" and smally = "0110011" else
			"111111" when smallx = "0010111" and smally = "0110011" else
			"111111" when smallx = "0011100" and smally = "0110011" else
			"111111" when smallx = "0100001" and smally = "0110011" else
			"111111" when smallx = "0101000" and smally = "0110011" else
			"111111" when smallx = "0101111" and smally = "0110011" else
			"111111" when smallx = "0110011" and smally = "0110011" else
			"111111" when smallx = "0110110" and smally = "0110011" else
			"111111" when smallx = "0111000" and smally = "0110011" else
			"111111" when smallx = "0111011" and smally = "0110011" else
			"111111" when smallx = "0111111" and smally = "0110011" else
			"111111" when smallx = "0001101" and smally = "0110100" else
			"111111" when smallx = "0001110" and smally = "0110100" else
			"111111" when smallx = "0001111" and smally = "0110100" else
			"111111" when smallx = "0010010" and smally = "0110100" else
			"111111" when smallx = "0010011" and smally = "0110100" else
			"111111" when smallx = "0010100" and smally = "0110100" else
			"111111" when smallx = "0010111" and smally = "0110100" else
			"111111" when smallx = "0011000" and smally = "0110100" else
			"111111" when smallx = "0011001" and smally = "0110100" else
			"111111" when smallx = "0011101" and smally = "0110100" else
			"111111" when smallx = "0011110" and smally = "0110100" else
			"111111" when smallx = "0100010" and smally = "0110100" else
			"111111" when smallx = "0100011" and smally = "0110100" else
			"111111" when smallx = "0101001" and smally = "0110100" else
			"111111" when smallx = "0101010" and smally = "0110100" else
			"111111" when smallx = "0101111" and smally = "0110100" else
			"111111" when smallx = "0110011" and smally = "0110100" else
			"111111" when smallx = "0110100" and smally = "0110100" else
			"111111" when smallx = "0110101" and smally = "0110100" else
			"111111" when smallx = "0110110" and smally = "0110100" else
			"111111" when smallx = "0111000" and smally = "0110100" else
			"111111" when smallx = "0111001" and smally = "0110100" else
			"111111" when smallx = "0111010" and smally = "0110100" else
			"111111" when smallx = "0111111" and smally = "0110100" else
			"111111" when smallx = "0001101" and smally = "0110101" else
			"111111" when smallx = "0010010" and smally = "0110101" else
			"111111" when smallx = "0010100" and smally = "0110101" else
			"111111" when smallx = "0010111" and smally = "0110101" else
			"111111" when smallx = "0011111" and smally = "0110101" else
			"111111" when smallx = "0100100" and smally = "0110101" else
			"111111" when smallx = "0101011" and smally = "0110101" else
			"111111" when smallx = "0101111" and smally = "0110101" else
			"111111" when smallx = "0110011" and smally = "0110101" else
			"111111" when smallx = "0110110" and smally = "0110101" else
			"111111" when smallx = "0111000" and smally = "0110101" else
			"111111" when smallx = "0111010" and smally = "0110101" else
			"111111" when smallx = "0111111" and smally = "0110101" else
			"111111" when smallx = "0001101" and smally = "0110110" else
			"111111" when smallx = "0010010" and smally = "0110110" else
			"111111" when smallx = "0010101" and smally = "0110110" else
			"111111" when smallx = "0010111" and smally = "0110110" else
			"111111" when smallx = "0011000" and smally = "0110110" else
			"111111" when smallx = "0011001" and smally = "0110110" else
			"111111" when smallx = "0011010" and smally = "0110110" else
			"111111" when smallx = "0011100" and smally = "0110110" else
			"111111" when smallx = "0011101" and smally = "0110110" else
			"111111" when smallx = "0011110" and smally = "0110110" else
			"111111" when smallx = "0100001" and smally = "0110110" else
			"111111" when smallx = "0100010" and smally = "0110110" else
			"111111" when smallx = "0100011" and smally = "0110110" else
			"111111" when smallx = "0101000" and smally = "0110110" else
			"111111" when smallx = "0101001" and smally = "0110110" else
			"111111" when smallx = "0101010" and smally = "0110110" else
			"111111" when smallx = "0101111" and smally = "0110110" else
			"111111" when smallx = "0110011" and smally = "0110110" else
			"111111" when smallx = "0110110" and smally = "0110110" else
			"111111" when smallx = "0111000" and smally = "0110110" else
			"111111" when smallx = "0111011" and smally = "0110110" else
			"111111" when smallx = "0111111" and smally = "0110110" else
			"011011";
end if;
end process;
end;
